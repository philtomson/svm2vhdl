--use std.textio.all;
--library ieee;
--use ieee.std_logic_1164.all;
--use work.numeric_std.all;


entity tb_csvm is
  generic(
    SV_ADDR_BITS     : natural := 9;
    SV_DATA_BITS     : natural := 18;
    SV_BINPT         : natural := 16; 

    XIN_ADDR_BITS    : natural := 1;
    XIN_DATA_BITS    : natural := 18;
    XIN_BINPT        : natural := 16;

    EXPLUT_ADDR_BITS : natural := 7;
    EXPLUT_DATA_BITS : natural := 16;
    EXPLUT_BINPT     : natural := 16;

    ALPHA_ADDR_BITS  : natural := 8;
    ALPHA_DATA_BITS  : natural := 17;
    ALPHA_BINPT      : natural := 16;

    RESULT_WIDTH     : natural := 33;

     

    DIFF_WIDTH       : natural := 18;
    
    DIFF_BINPT       : natural := 16;
    
    DIFF_SQUARED_WIDTH : natural := 36;
    
    DIFF_SQUARED_BINPT: natural := 32;
    
    --KWIDTH           : natural := 35;
    --KBINPT           : natural := 32;
    KWIDTH           : natural := 18;
    KBINPT           : natural := 16;
    
    EXPXALPHA_BITS   : natural := 33;
    EXPXALPHA_BINPT  : natural := 32;
    ACCUM_BITS       : natural := 40;
    ACCUM_BINPT      : natural := 16;

    NSV              : natural := 242;
    NI               : natural := 2  );
end tb_csvm;

use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


----------------------------------------------------------------
-- xin values:
-- 0:xin(0): 0.86195129   "00.1101110010101001"
-- 0:xin(1): -1.2353323   "10.1100001111000001"
----------------------------------------------------------------
-- 1:xin(0): 0.90818191   "00.1110100001111111"    
-- 1:xin(1): 1.4833819    "01.0111101110111111"
----------------------------------------------------------------
-- 2:xin(0): 0.07448764   "00.0001001100010010"  
-- 2:xin(1): -0.60681143  "11.0110010010101000
----------------------------------------------------------------
-- 3:xin(0): 0.735740819074673 "00.1011110001011010" 
-- 3:xin(1): 0.475955584677872 "00.0111100111011000"

architecture testbench of tb_csvm is

type test_vector is record
  xin_0: signed(XIN_DATA_BITS -1 downto 0); xin_1: signed(XIN_DATA_BITS -1 downto 0); pass: boolean;
end record;
type test_vector_array is array(natural range <>) of test_vector;
constant test_vectors: test_vector_array := (
--  (xin_0 => "001011011100110110", xin_1 => "000010011110001111", pass => true),
--  (xin_0 => "001001001010110100", xin_1 => "000100011000100000", pass => true),
--  (xin_0 => "001011110001011010", xin_1 => "000111100111011000", pass => false),
  (xin_0 => "000010110010110110", xin_1 => "000000100110011100", pass => true),
  (xin_0 => "001000111000100111", xin_1 => "000011001011101110", pass => false),
  (xin_0 => "000111100100110011", xin_1 => "000001101011111011", pass => false),
  (xin_0 => "000100010001010010", xin_1 => "001000000010000001", pass => false),
  (xin_0 => "000101001110100111", xin_1 => "000101011011010010", pass => true),
  (xin_0 => "001001010111100110", xin_1 => "001001011011010101", pass => false),
  (xin_0 => "001010110110110000", xin_1 => "001000110010110011", pass => false),
  (xin_0 => "000111010101010110", xin_1 => "000110011010001000", pass => true),
  (xin_0 => "001100100101111011", xin_1 => "001000101001111110", pass => false),
  (xin_0 => "001110011000101000", xin_1 => "001001110101010010", pass => true),
  (xin_0 => "001000001010101100", xin_1 => "001011000011101000", pass => false),
  (xin_0 => "001000010101000101", xin_1 => "000111111001010111", pass => true),
  (xin_0 => "001010001010001110", xin_1 => "000110100010000111", pass => true),
  (xin_0 => "000100000111110011", xin_1 => "000000111101100101", pass => true),
  (xin_0 => "001010010010111110", xin_1 => "000011110100100101", pass => true),
  (xin_0 => "000111010011101001", xin_1 => "000010000101011110", pass => false),
  (xin_0 => "000110110010001010", xin_1 => "001010000010110010", pass => false),
  (xin_0 => "001010111010101001", xin_1 => "001001001010001000", pass => false),
  (xin_0 => "001001011101100110", xin_1 => "001001111101111010", pass => false),
  (xin_0 => "001100100010000100", xin_1 => "001000111111001100", pass => false),
  (xin_0 => "000110000010001100", xin_1 => "000101000001010111", pass => true),
  (xin_0 => "000110101000000000", xin_1 => "000011110110011000", pass => false),
  (xin_0 => "001000011110000111", xin_1 => "001001011110100010", pass => false),
  (xin_0 => "001101111000101001", xin_1 => "000100100010101101", pass => false),
  (xin_0 => "001000011100101010", xin_1 => "000100110001100100", pass => true),
  (xin_0 => "001001111011111111", xin_1 => "000011000111000000", pass => false),
  (xin_0 => "001010000111001011", xin_1 => "000001111111011100", pass => false),
  (xin_0 => "001100111101001101", xin_1 => "000101011111000011", pass => false),
  (xin_0 => "001100000101100110", xin_1 => "001000101000010010", pass => false),
  (xin_0 => "000110000111111010", xin_1 => "001000001010110100", pass => true),
  (xin_0 => "001000110101010000", xin_1 => "000011000111001010", pass => false),
  (xin_0 => "001010100100010110", xin_1 => "000011000100111011", pass => true),
  (xin_0 => "000010101000100001", xin_1 => "000000100001011101", pass => true),
  (xin_0 => "000101010111111100", xin_1 => "000111001101011110", pass => true),
  (xin_0 => "000101110100010000", xin_1 => "000111010011111010", pass => true),
  (xin_0 => "000111100101011001", xin_1 => "000110001010101101", pass => true),
  (xin_0 => "001011001101010110", xin_1 => "001001000111101100", pass => false),
  (xin_0 => "000110011101011100", xin_1 => "000010011000010011", pass => false),
  (xin_0 => "000110110011110001", xin_1 => "000001100101110101", pass => false),
  (xin_0 => "000101011100001001", xin_1 => "000111010100000011", pass => true),
  (xin_0 => "001011011010000010", xin_1 => "000100010111111101", pass => true),
  (xin_0 => "001001010001000010", xin_1 => "000101010011011000", pass => true),
  (xin_0 => "001011011001001000", xin_1 => "000101000110001110", pass => true),
  (xin_0 => "001000111000000011", xin_1 => "000010111001110110", pass => false),
  (xin_0 => "000110011111001101", xin_1 => "000110110011010100", pass => true),
  (xin_0 => "000110001100100110", xin_1 => "001010011101000010", pass => false),
  (xin_0 => "000110111000010001", xin_1 => "000101101000111010", pass => true),
  (xin_0 => "000011010000001101", xin_1 => "001000000101100000", pass => false),
  (xin_0 => "001011011000110111", xin_1 => "000101101100011011", pass => true),
  (xin_0 => "001010001001010001", xin_1 => "001010101011110111", pass => false),
  (xin_0 => "000101111101100000", xin_1 => "001000001101111000", pass => false),
  (xin_0 => "001100010001101001", xin_1 => "000001011111001001", pass => true),
  (xin_0 => "001000010110111000", xin_1 => "000010101110001111", pass => false),
  (xin_0 => "000111010110001001", xin_1 => "001000111111010001", pass => false),
  (xin_0 => "000100101011110101", xin_1 => "000111110011110011", pass => false),
  (xin_0 => "001101111000001001", xin_1 => "000110001000000010", pass => false),
  (xin_0 => "000101011101011101", xin_1 => "001001010001100011", pass => false),
  (xin_0 => "000110100101111010", xin_1 => "000100001001111100", pass => true),
  (xin_0 => "000101110100100000", xin_1 => "000011010101010100", pass => false),
  (xin_0 => "001100101010110011", xin_1 => "000101100000101011", pass => false),
  (xin_0 => "000111011000011111", xin_1 => "001001101000000001", pass => false),
  (xin_0 => "001000001100000010", xin_1 => "000110011001101010", pass => true),
  (xin_0 => "000101100100110100", xin_1 => "000011010101101010", pass => true),
  (xin_0 => "001000000000100010", xin_1 => "000110011101100001", pass => true),
  (xin_0 => "001010110101000001", xin_1 => "000111001100001011", pass => false),
  (xin_0 => "000011101101110011", xin_1 => "000100101111101100", pass => true),
  (xin_0 => "000111100000000010", xin_1 => "001001100011100110", pass => false),
  (xin_0 => "000010100111000111", xin_1 => "000110100001110110", pass => false),
  (xin_0 => "001000011100100000", xin_1 => "000110011011000110", pass => true),
  (xin_0 => "001010010100100011", xin_1 => "000110100001100111", pass => true),
  (xin_0 => "000111111000100000", xin_1 => "000011001111001011", pass => false),
  (xin_0 => "001011001100100011", xin_1 => "000010100001001000", pass => true),
  (xin_0 => "001001010101110000", xin_1 => "001100011101000001", pass => false),
  (xin_0 => "001000100111111101", xin_1 => "001000110011000111", pass => true),
  (xin_0 => "001000010000101110", xin_1 => "000001111011001110", pass => false),
  (xin_0 => "001010011100110111", xin_1 => "001011011011111011", pass => false),
  (xin_0 => "001011100111011011", xin_1 => "001000101001101110", pass => false),
  (xin_0 => "000101111101001100", xin_1 => "000111000100011110", pass => true),
  (xin_0 => "001010101000011110", xin_1 => "001001110001011001", pass => false),
  (xin_0 => "000101011001011111", xin_1 => "000101010010100111", pass => true),
  (xin_0 => "001010100011101010", xin_1 => "000100110110001101", pass => true),
  (xin_0 => "001011101010000100", xin_1 => "001000011000111011", pass => false),
  (xin_0 => "001011110110110011", xin_1 => "000110111111111110", pass => false),
  (xin_0 => "001100110101010101", xin_1 => "000110100001111110", pass => false),
  (xin_0 => "000110110011100001", xin_1 => "001001001101000011", pass => false),
  (xin_0 => "000111101001010011", xin_1 => "001000011011001100", pass => true),
  (xin_0 => "000100001100010101", xin_1 => "000110101010011000", pass => true),
  (xin_0 => "001001001110111110", xin_1 => "001000000001001001", pass => true),
  (xin_0 => "001001001111000011", xin_1 => "000010001011110110", pass => false),
  (xin_0 => "000101111000100000", xin_1 => "000001100010011011", pass => false),
  (xin_0 => "001101001000010001", xin_1 => "000111010100001010", pass => false),
  (xin_0 => "001001000110110011", xin_1 => "001010110110010111", pass => false),
  (xin_0 => "001010110011000111", xin_1 => "001001001110000010", pass => false),
  (xin_0 => "001101001011000110", xin_1 => "001011010110100010", pass => true),
  (xin_0 => "001000101000101100", xin_1 => "000011011101010010", pass => false),
  (xin_0 => "001100000110100100", xin_1 => "000111001000101110", pass => false),
  (xin_0 => "001001111100111011", xin_1 => "000011100001001101", pass => false),
  (xin_0 => "001110100111010001", xin_1 => "001000111110000100", pass => true),
  (xin_0 => "001001000010100000", xin_1 => "001001111000001010", pass => false),
  (xin_0 => "001011011111011100", xin_1 => "000011110001011110", pass => true),
  (xin_0 => "001000010011000101", xin_1 => "000001110011101101", pass => false),
  (xin_0 => "001001000011010000", xin_1 => "000010110010101010", pass => false),
  (xin_0 => "001010101000010100", xin_1 => "000011000111100100", pass => true),
  (xin_0 => "001001001001001111", xin_1 => "000010011111111000", pass => false),
  (xin_0 => "001011011001011110", xin_1 => "000101000000010001", pass => true),
  (xin_0 => "000111110010110110", xin_1 => "000010000100111100", pass => false),
  (xin_0 => "001010001001101110", xin_1 => "001001101111101111", pass => false),
  (xin_0 => "000011110100110001", xin_1 => "000011101101011010", pass => true),
  (xin_0 => "001011000011011010", xin_1 => "000100100101100001", pass => true),
  (xin_0 => "000111001010010101", xin_1 => "000010100110000001", pass => false),
  (xin_0 => "001000111000101100", xin_1 => "000010011110000100", pass => false),
  (xin_0 => "001000110011001010", xin_1 => "000010011001010011", pass => false),
  (xin_0 => "001101000110111001", xin_1 => "000010100100000101", pass => true),
  (xin_0 => "001000111011111001", xin_1 => "000101010000010101", pass => true),
  (xin_0 => "000111000110100110", xin_1 => "001010001111000111", pass => false),
  (xin_0 => "001010011010011100", xin_1 => "001011101000011001", pass => false),
  (xin_0 => "000100011100100011", xin_1 => "000010111001001111", pass => true),
  (xin_0 => "001100001110000110", xin_1 => "000110001100010011", pass => false),
  (xin_0 => "000111010111111000", xin_1 => "000010001110111110", pass => false),
  (xin_0 => "000101100100011110", xin_1 => "000110111001101011", pass => true),
  (xin_0 => "001100111100101100", xin_1 => "000110101000000111", pass => false),
  (xin_0 => "001100011010011101", xin_1 => "001000010110001010", pass => false),
  (xin_0 => "000101110100111111", xin_1 => "001001010011100110", pass => false),
  (xin_0 => "001100011101011010", xin_1 => "000110110100111101", pass => false),
  (xin_0 => "001000101100101001", xin_1 => "001001110001101001", pass => false),
  (xin_0 => "000111011110100011", xin_1 => "000011011001001101", pass => false),
  (xin_0 => "000111101010010100", xin_1 => "000010010110011010", pass => false),
  (xin_0 => "001001001111100011", xin_1 => "000001101111000001", pass => false),
  (xin_0 => "001000001010111111", xin_1 => "000010010100110110", pass => false),
  (xin_0 => "000111011010111101", xin_1 => "000011000111010001", pass => false),
  (xin_0 => "000110001110000100", xin_1 => "000010011001101010", pass => false),
  (xin_0 => "000110101011001110", xin_1 => "000011001000000110", pass => false),
  (xin_0 => "001010001100111011", xin_1 => "000010001100000001", pass => false),
  (xin_0 => "001000000101010011", xin_1 => "000011000100111101", pass => false),
  (xin_0 => "001000001110011110", xin_1 => "000111001110001000", pass => true),
  (xin_0 => "001100000010111101", xin_1 => "000101100011100011", pass => true),
  (xin_0 => "001010101110011110", xin_1 => "001010011001101101", pass => false),
  (xin_0 => "000111100001000001", xin_1 => "001010100000001010", pass => false),
  (xin_0 => "001010100011010010", xin_1 => "001100011101001010", pass => false),
  (xin_0 => "001000010001011111", xin_1 => "000111010010111101", pass => true),
  (xin_0 => "001101110111110111", xin_1 => "001001111001001101", pass => true),
  (xin_0 => "001100010111110001", xin_1 => "000111001111011101", pass => false),
  (xin_0 => "001011011010110001", xin_1 => "001010101011100001", pass => false),
  (xin_0 => "001100001001010101", xin_1 => "000101000101101111", pass => true),
  (xin_0 => "001000101000110010", xin_1 => "000010111110111100", pass => false),
  (xin_0 => "000010011011011011", xin_1 => "000000010000101011", pass => true),
  (xin_0 => "000101111101101101", xin_1 => "001001110100011010", pass => false),
  (xin_0 => "000110010001101000", xin_1 => "001010101001010110", pass => false),
  (xin_0 => "000111010100000001", xin_1 => "001001110101100110", pass => false),
  (xin_0 => "001011011110001000", xin_1 => "000111111110100101", pass => false),
  (xin_0 => "001100111110110011", xin_1 => "000111000001100010", pass => false),
  (xin_0 => "001011000110001001", xin_1 => "001100101110010111", pass => false),
  (xin_0 => "001101000011100100", xin_1 => "000101110010001111", pass => false),
  (xin_0 => "000111011100100101", xin_1 => "000010101011110010", pass => false),
  (xin_0 => "001011101000001111", xin_1 => "000011001000101000", pass => true),
  (xin_0 => "000101111110000111", xin_1 => "001000010010111111", pass => false),
  (xin_0 => "001111111001111111", xin_1 => "001001110111010111", pass => true),
  (xin_0 => "000011001101101111", xin_1 => "001000111000110100", pass => false),
  (xin_0 => "000011111010001011", xin_1 => "000000101010000001", pass => true),
  (xin_0 => "001010011110001011", xin_1 => "000101100001101100", pass => true),
  (xin_0 => "001001000011011011", xin_1 => "001011011001001010", pass => false),
  (xin_0 => "001001110111011100", xin_1 => "000101101011001001", pass => true),
  (xin_0 => "001010001110100111", xin_1 => "001000111101101101", pass => false),
  (xin_0 => "001101010001001010", xin_1 => "001010111011010011", pass => true),
  (xin_0 => "001011100101100111", xin_1 => "000110100101011111", pass => false),
  (xin_0 => "001000011011110100", xin_1 => "000110110011011110", pass => true),
  (xin_0 => "001100110000000101", xin_1 => "000111001110010101", pass => false),
  (xin_0 => "001010100101111100", xin_1 => "000110011110011011", pass => true),
  (xin_0 => "000100101000000001", xin_1 => "000110001001011001", pass => true),
  (xin_0 => "001101010101010000", xin_1 => "001011000011111001", pass => true),
  (xin_0 => "001001110101010011", xin_1 => "000110001101110011", pass => true),
  (xin_0 => "000110001010101101", xin_1 => "000101111010101110", pass => true),
  (xin_0 => "000111100010000101", xin_1 => "000001110011110111", pass => false),
  (xin_0 => "000111100001001101", xin_1 => "001010001101000110", pass => false),
  (xin_0 => "001001111110100100", xin_1 => "001001011101011001", pass => false),
  (xin_0 => "000100111011101001", xin_1 => "000101110000010011", pass => true),
  (xin_0 => "001100111010001000", xin_1 => "000111101100011001", pass => false),
  (xin_0 => "001010101011001101", xin_1 => "001011101101011011", pass => false),
  (xin_0 => "001000010010010010", xin_1 => "000011001001000001", pass => false),
  (xin_0 => "001000110101110011", xin_1 => "000011001111000101", pass => false),
  (xin_0 => "001001110011000101", xin_1 => "000101101111101110", pass => true),
  (xin_0 => "001011110110101111", xin_1 => "001000001101101110", pass => false),
  (xin_0 => "001000100101111100", xin_1 => "000110110001110101", pass => true),
  (xin_0 => "001001010001111101", xin_1 => "000111101000011000", pass => true),
  (xin_0 => "000110011111010011", xin_1 => "000011011011100101", pass => false),
  (xin_0 => "000100111011001000", xin_1 => "000101110111100001", pass => true),
  (xin_0 => "000100101101100110", xin_1 => "001000000010000011", pass => false),
  (xin_0 => "001110001010011001", xin_1 => "000110011010011000", pass => false),
  (xin_0 => "001010000000100010", xin_1 => "000011100111101001", pass => false),
  (xin_0 => "000111100000111011", xin_1 => "001001011110000101", pass => false),
  (xin_0 => "000011101001100111", xin_1 => "000011010010111110", pass => true),
  (xin_0 => "000110111110011011", xin_1 => "000110101001101100", pass => true),
  (xin_0 => "001011110111110001", xin_1 => "001000110110110011", pass => false),
  (xin_0 => "000011101110101001", xin_1 => "000001010010100011", pass => true),
  (xin_0 => "000100111111001000", xin_1 => "000101101100000011", pass => true),
  (xin_0 => "001100011011110011", xin_1 => "000100001010010100", pass => true),
  (xin_0 => "001000001001010011", xin_1 => "000010011100000011", pass => false),
  (xin_0 => "000111011111111011", xin_1 => "000011000011111110", pass => false),
  (xin_0 => "001000110010111001", xin_1 => "000001110100000100", pass => false),
  (xin_0 => "001011000110101110", xin_1 => "000010101000001101", pass => true),
  (xin_0 => "001011100110110110", xin_1 => "001011001011101101", pass => false),
  (xin_0 => "001001010100100001", xin_1 => "001100000111111000", pass => false),
  (xin_0 => "001100000000010101", xin_1 => "001000100101100000", pass => false),
  (xin_0 => "000011110101100010", xin_1 => "000111100111100001", pass => false),
  (xin_0 => "000110011100111011", xin_1 => "000110110000011101", pass => true),
  (xin_0 => "000100101010001111", xin_1 => "001001000110001000", pass => false),
  (xin_0 => "000100111010011000", xin_1 => "000101001111111100", pass => true),
  (xin_0 => "001001101110101110", xin_1 => "001001101011111011", pass => false),
  (xin_0 => "000100011000010000", xin_1 => "000011110011010010", pass => true),
  (xin_0 => "001010101110101110", xin_1 => "001010010101100101", pass => false),
  (xin_0 => "001100011001010100", xin_1 => "000011010010101000", pass => true),
  (xin_0 => "000111000110100101", xin_1 => "001010000010011100", pass => false),
  (xin_0 => "001001011110111111", xin_1 => "000010101100001100", pass => false),
  (xin_0 => "001101000111111101", xin_1 => "000001000011100100", pass => true),
  (xin_0 => "000110110011000000", xin_1 => "000001111111110000", pass => false),
  (xin_0 => "000110101111110101", xin_1 => "000001110110000101", pass => false),
  (xin_0 => "001001010110000111", xin_1 => "000110011000111010", pass => true),
  (xin_0 => "000100111100011110", xin_1 => "000010110111011001", pass => true),
  (xin_0 => "001100101000001000", xin_1 => "000101101000101111", pass => false),
  (xin_0 => "001001000101000101", xin_1 => "000110010001000001", pass => true),
  (xin_0 => "000100111001011100", xin_1 => "000001100011010100", pass => true),
  (xin_0 => "000110100100010010", xin_1 => "001001100100101111", pass => false),
  (xin_0 => "001100101100111011", xin_1 => "000110101100010110", pass => false),
  (xin_0 => "001000111010111010", xin_1 => "000011110110110111", pass => false),
  (xin_0 => "001010101011111100", xin_1 => "000110101000010111", pass => true),
  (xin_0 => "000111001000000101", xin_1 => "001001000111001010", pass => false),
  (xin_0 => "000101001000101101", xin_1 => "000110010110010101", pass => true),
  (xin_0 => "001100010011011100", xin_1 => "000110011000000100", pass => false),
  (xin_0 => "001000100010001001", xin_1 => "001011001111010100", pass => false),
  (xin_0 => "001001001110111000", xin_1 => "000010000010100000", pass => false),
  (xin_0 => "000010111000110010", xin_1 => "000010100000110100", pass => true),
  (xin_0 => "001000111000011011", xin_1 => "000011111001101011", pass => false),
  (xin_0 => "001001100011010100", xin_1 => "001000001101000010", pass => true),
  (xin_0 => "001101001011010000", xin_1 => "000101110011011011", pass => false),
  (xin_0 => "001010010100110011", xin_1 => "000111010000011100", pass => true),
  (xin_0 => "001001001101010100", xin_1 => "000010011010111100", pass => false),
  (xin_0 => "001011111110110100", xin_1 => "000011010011111000", pass => true),
  (xin_0 => "001010100100111011", xin_1 => "000111101110000010", pass => false),
  (xin_0 => "000111001001110010", xin_1 => "001001100101101010", pass => false),
  (xin_0 => "001000010100100100", xin_1 => "000011000010011011", pass => false),
  (xin_0 => "001010000111000010", xin_1 => "000100011011000001", pass => true),
  (xin_0 => "001011100110110000", xin_1 => "000010010110101110", pass => true),
  (xin_0 => "001111000100100010", xin_1 => "001001000101110011", pass => true),
  (xin_0 => "001000010101110010", xin_1 => "000101110000011100", pass => true),
  (xin_0 => "000110100111100011", xin_1 => "000111111110011000", pass => true),
  (xin_0 => "001010110011001100", xin_1 => "000110001111100111", pass => true),
  (xin_0 => "001000111011110101", xin_1 => "000011001011101111", pass => false),
  (xin_0 => "001010010101100010", xin_1 => "000010011101111111", pass => false),
  (xin_0 => "001010101111000000", xin_1 => "000111010111100111", pass => false),
  (xin_0 => "001101001100000011", xin_1 => "000010001110000100", pass => true),
  (xin_0 => "001100001101000110", xin_1 => "001000000101100011", pass => false),
  (xin_0 => "000100010100000100", xin_1 => "001000010011010010", pass => false),
  (xin_0 => "000101000110000000", xin_1 => "001000011010011011", pass => false),
  (xin_0 => "001110101101000100", xin_1 => "000110001001101010", pass => false),
  (xin_0 => "000111011111101100", xin_1 => "001010010101111100", pass => false),
  (xin_0 => "001010010100001111", xin_1 => "001001111001111010", pass => false),
  (xin_0 => "001111010101100110", xin_1 => "001001101100001010", pass => true),
  (xin_0 => "000111110011010000", xin_1 => "000010010110000001", pass => false),
  (xin_0 => "000011110101010111", xin_1 => "000100110110000011", pass => true),
  (xin_0 => "001011110001111001", xin_1 => "000010001001000001", pass => true),
  (xin_0 => "001010000101010000", xin_1 => "001010000100110000", pass => false),
  (xin_0 => "001100100110110001", xin_1 => "000101001110101111", pass => true),
  (xin_0 => "000111111000000001", xin_1 => "001010111010100000", pass => false),
  (xin_0 => "000101011110100001", xin_1 => "000011101101111101", pass => true),
  (xin_0 => "000000010100001110", xin_1 => "000101101111100001", pass => false),
  (xin_0 => "000111001101100110", xin_1 => "000100100101100111", pass => true),
  (xin_0 => "001001100001011011", xin_1 => "001011100100111010", pass => false),
  (xin_0 => "000011010110100111", xin_1 => "000011011011100000", pass => true),
  (xin_0 => "000110000001100100", xin_1 => "000010011110101010", pass => false),
  (xin_0 => "000110101001101011", xin_1 => "001001011110101011", pass => false),
  (xin_0 => "000111010001011001", xin_1 => "000100011101111010", pass => true),
  (xin_0 => "000111000001000101", xin_1 => "001001000001011010", pass => false),
  (xin_0 => "000110110001011100", xin_1 => "000110000010100111", pass => true),
  (xin_0 => "000110110100100110", xin_1 => "001000010011011011", pass => true),
  (xin_0 => "001011100000101011", xin_1 => "001000000010111000", pass => false),
  (xin_0 => "000011010110110001", xin_1 => "001000000011111010", pass => false),
  (xin_0 => "001100011101101000", xin_1 => "000110011000100001", pass => false),
  (xin_0 => "000100111010010111", xin_1 => "001001100011011011", pass => false),
  (xin_0 => "000101010010101110", xin_1 => "000101110111010100", pass => true),
  (xin_0 => "001010101101110110", xin_1 => "000110010001001011", pass => true),
  (xin_0 => "001101001010101011", xin_1 => "000000110101001000", pass => true),
  (xin_0 => "000100010010111100", xin_1 => "000101001000000001", pass => true),
  (xin_0 => "000110000011001110", xin_1 => "000110011101110000", pass => true),
  (xin_0 => "000111011001101100", xin_1 => "001001110110111001", pass => false),
  (xin_0 => "000011111100011101", xin_1 => "001000110111111010", pass => false),
  (xin_0 => "000100000111110000", xin_1 => "000101100101010011", pass => true),
  (xin_0 => "000101111011101101", xin_1 => "001000010010101100", pass => false),
  (xin_0 => "001101100111101111", xin_1 => "000101000011010011", pass => false),
  (xin_0 => "001100001111010111", xin_1 => "000010010111110001", pass => true),
  (xin_0 => "001100011101100101", xin_1 => "000011001000000000", pass => true),
  (xin_0 => "001011110001100100", xin_1 => "000001110000011001", pass => true),
  (xin_0 => "001001010011000011", xin_1 => "000010010101100111", pass => false),
  (xin_0 => "001100001010001111", xin_1 => "001000010011101111", pass => false),
  (xin_0 => "001001111001101110", xin_1 => "000110101111101101", pass => true),
  (xin_0 => "001011110011011000", xin_1 => "000110110101111111", pass => false),
  (xin_0 => "001010000111011001", xin_1 => "000010001111000111", pass => false),
  (xin_0 => "001100011100010111", xin_1 => "000001011110110011", pass => true),
  (xin_0 => "000100011101001111", xin_1 => "000111011000001100", pass => false),
  (xin_0 => "000100100100110010", xin_1 => "000101101000010110", pass => true),
  (xin_0 => "000110010010110011", xin_1 => "001010100110100111", pass => false),
  (xin_0 => "001001101111111111", xin_1 => "001001110011011100", pass => false),
  (xin_0 => "001001100011100000", xin_1 => "000010100010110011", pass => false),
  (xin_0 => "001011111010101111", xin_1 => "000110100001100010", pass => false),
  (xin_0 => "001000111011000001", xin_1 => "000011010011101101", pass => false),
  (xin_0 => "001100000010011111", xin_1 => "000100111011011001", pass => true),
  (xin_0 => "000011011110010111", xin_1 => "000001000100100111", pass => true),
  (xin_0 => "001111101111011110", xin_1 => "001001101010001110", pass => true),
  (xin_0 => "001100101110001101", xin_1 => "001000011110011001", pass => false),
  (xin_0 => "000110001100110101", xin_1 => "000110101010011111", pass => true),
  (xin_0 => "000111101010010110", xin_1 => "000001100101000101", pass => false),
  (xin_0 => "000100110011001111", xin_1 => "000100100100010110", pass => true),
  (xin_0 => "001100101110111000", xin_1 => "000110110000101100", pass => false),
  (xin_0 => "001000100101001001", xin_1 => "001010111111110010", pass => false),
  (xin_0 => "001010111111010101", xin_1 => "000100011101001010", pass => true),
  (xin_0 => "001011111010001001", xin_1 => "001000011010101010", pass => false),
  (xin_0 => "000011011111000100", xin_1 => "000100111101010101", pass => true),
  (xin_0 => "000110000100100011", xin_1 => "000011101100101001", pass => false),
  (xin_0 => "000100101101011111", xin_1 => "001001100110111110", pass => false),
  (xin_0 => "001011111100110011", xin_1 => "001000101011010000", pass => false),
  (xin_0 => "001100111110010111", xin_1 => "000110011010011010", pass => false),
  (xin_0 => "001010101011010001", xin_1 => "001000010010010010", pass => false),
  (xin_0 => "001001011001110101", xin_1 => "001011111011101010", pass => false),
  (xin_0 => "001001110001100010", xin_1 => "000001011111001101", pass => false),
  (xin_0 => "001001100010011000", xin_1 => "000010000011001111", pass => false),
  (xin_0 => "001011001001010111", xin_1 => "000101100110000100", pass => true),
  (xin_0 => "001001010101100100", xin_1 => "000001101100111100", pass => false),
  (xin_0 => "001011101001001110", xin_1 => "000011011111000010", pass => true),
  (xin_0 => "000110111110110010", xin_1 => "000100011100100011", pass => true),
  (xin_0 => "000101100010100000", xin_1 => "000110010100011100", pass => true),
  (xin_0 => "001100011001100100", xin_1 => "000010001010011010", pass => true),
  (xin_0 => "000110011101111001", xin_1 => "000010100101100101", pass => false),
  (xin_0 => "001110011010100001", xin_1 => "000111001101101110", pass => false),
  (xin_0 => "001000000010101110", xin_1 => "000011011011110111", pass => false),
  (xin_0 => "000110110111000011", xin_1 => "001001110110000110", pass => false),
  (xin_0 => "000010110000000100", xin_1 => "000001011001111000", pass => true),
  (xin_0 => "000111011001001001", xin_1 => "000010101110110010", pass => false),
  (xin_0 => "001000010110010110", xin_1 => "000111001111001010", pass => true),
  (xin_0 => "001010001111111011", xin_1 => "001001000001011111", pass => false),
  (xin_0 => "000100100010110011", xin_1 => "000110001101111010", pass => true),
  (xin_0 => "000100011001000010", xin_1 => "001000111110101101", pass => false),
  (xin_0 => "000110101110010001", xin_1 => "000111010101011011", pass => true),
  (xin_0 => "001100100111111101", xin_1 => "000111001001001010", pass => false),
  (xin_0 => "001000101101010101", xin_1 => "001001101110001101", pass => false),
  (xin_0 => "000111101110011010", xin_1 => "000110010010100101", pass => true),
  (xin_0 => "000101100010010111", xin_1 => "001000011101000001", pass => false),
  (xin_0 => "000110001011010110", xin_1 => "001000101100100011", pass => false),
  (xin_0 => "001000101110100000", xin_1 => "000010111001011011", pass => false),
  (xin_0 => "000011101000100010", xin_1 => "000011101010000000", pass => true),
  (xin_0 => "000111111111001000", xin_1 => "000010001010001111", pass => false),
  (xin_0 => "000111100001111000", xin_1 => "000001100000100101", pass => false),
  (xin_0 => "001011010001010101", xin_1 => "001010111110111011", pass => false),
  (xin_0 => "001110000001101011", xin_1 => "001010010001110111", pass => true),
  (xin_0 => "001010110111100110", xin_1 => "001011011000000010", pass => false),
  (xin_0 => "000111110011111000", xin_1 => "000101011101010000", pass => true),
  (xin_0 => "000101010111001011", xin_1 => "001000100111110111", pass => false),
  (xin_0 => "000111100101010010", xin_1 => "000011111100110001", pass => false),
  (xin_0 => "001001111011111011", xin_1 => "001000111001111010", pass => false),
  (xin_0 => "001100001110111111", xin_1 => "000111001110110100", pass => false),
  (xin_0 => "000111011010101010", xin_1 => "000011010110111000", pass => false),
  (xin_0 => "000101100101001000", xin_1 => "001001010110000101", pass => false),
  (xin_0 => "001000100011001110", xin_1 => "000110101000010101", pass => true),
  (xin_0 => "001000111101100001", xin_1 => "000011010001010001", pass => false),
  (xin_0 => "001011101011100101", xin_1 => "001010101010010110", pass => false),
  (xin_0 => "001100100010011111", xin_1 => "000100001000110111", pass => true),
  (xin_0 => "001100001010111100", xin_1 => "000100110001111001", pass => true),
  (xin_0 => "001000001100011101", xin_1 => "000010100101101101", pass => false),
  (xin_0 => "000111111101011000", xin_1 => "000001111111111011", pass => false),
  (xin_0 => "001011010100111101", xin_1 => "000110010111100100", pass => true),
  (xin_0 => "001010010011011000", xin_1 => "000111001101001111", pass => true),
  (xin_0 => "001001100010010011", xin_1 => "000110001111000010", pass => true),
  (xin_0 => "000100100110011010", xin_1 => "000010100000100001", pass => true),
  (xin_0 => "001001010100011100", xin_1 => "000010111100011001", pass => false),
  (xin_0 => "001000000111100101", xin_1 => "000111001001111001", pass => true),
  (xin_0 => "001011110011101010", xin_1 => "001001110000010001", pass => false),
  (xin_0 => "001001110100011011", xin_1 => "000011101111001001", pass => false),
  (xin_0 => "001011010011111011", xin_1 => "001000101101011110", pass => false),
  (xin_0 => "000111000110011101", xin_1 => "001000010010110101", pass => true),
  (xin_0 => "001000111100101100", xin_1 => "000111000101011011", pass => true),
  (xin_0 => "001000100110011110", xin_1 => "000110000001100000", pass => true),
  (xin_0 => "000110011100010000", xin_1 => "000110111000001100", pass => true),
  (xin_0 => "001111100001111101", xin_1 => "000111000101110100", pass => false),
  (xin_0 => "001001101001110111", xin_1 => "000111010010000100", pass => true),
  (xin_0 => "001011010001001110", xin_1 => "000011001110000001", pass => true),
  (xin_0 => "001000110001010000", xin_1 => "000100000110100100", pass => false),
  (xin_0 => "000110011101001010", xin_1 => "001010110111011111", pass => false),
  (xin_0 => "001100101111011101", xin_1 => "000101011101001010", pass => false),
  (xin_0 => "001001111001010110", xin_1 => "000110001000001111", pass => true),
  (xin_0 => "000111110101010101", xin_1 => "000111000001001110", pass => true),
  (xin_0 => "001100011101101001", xin_1 => "001000001011011111", pass => false),
  (xin_0 => "001000111001100000", xin_1 => "000010010101011000", pass => false),
  (xin_0 => "001011010001100101", xin_1 => "001001101011100100", pass => false),
  (xin_0 => "000011100001011000", xin_1 => "000111010111001010", pass => false),
  (xin_0 => "001000111111001000", xin_1 => "001011010001101000", pass => false),
  (xin_0 => "001010101000001010", xin_1 => "000100010101100100", pass => true),
  (xin_0 => "001000111011110110", xin_1 => "000011010011111011", pass => false),
  (xin_0 => "001011101010000100", xin_1 => "001000011001111101", pass => false),
  (xin_0 => "000100011010000111", xin_1 => "000101000000100100", pass => true),
  (xin_0 => "000100110000010011", xin_1 => "000110000101100101", pass => true),
  (xin_0 => "001100001011101111", xin_1 => "000101111010000001", pass => false),
  (xin_0 => "001001111100110111", xin_1 => "001010110000011011", pass => false),
  (xin_0 => "001000111111110111", xin_1 => "000001111101000011", pass => false),
  (xin_0 => "000101000111010010", xin_1 => "000101110111001100", pass => true),
  (xin_0 => "001011001110010101", xin_1 => "001010011100100110", pass => false),
  (xin_0 => "000110101000101100", xin_1 => "001011010000111010", pass => false),
  (xin_0 => "000101010011010100", xin_1 => "000011001010010001", pass => true),
  (xin_0 => "001101111001011001", xin_1 => "001001110010011111", pass => true),
  (xin_0 => "001001000001000100", xin_1 => "000101000011000111", pass => true),
  (xin_0 => "001000101111001101", xin_1 => "000100110100100011", pass => true),
  (xin_0 => "001000110011001100", xin_1 => "000110001011010011", pass => true),
  (xin_0 => "010000000000001100", xin_1 => "001010011101110111", pass => true),
  (xin_0 => "000100001000011000", xin_1 => "000100100001100100", pass => true),
  (xin_0 => "000110010010001110", xin_1 => "000010100111011010", pass => false),
  (xin_0 => "001001010001110010", xin_1 => "000110111100111011", pass => true),
  (xin_0 => "000110111111001111", xin_1 => "000100111101011110", pass => true),
  (xin_0 => "000100100000001010", xin_1 => "001000010011110011", pass => false),
  (xin_0 => "000101110100000110", xin_1 => "000110000011000000", pass => true),
  (xin_0 => "001100010001011110", xin_1 => "000111001110100111", pass => false),
  (xin_0 => "000101001001100100", xin_1 => "000110111101000111", pass => true),
  (xin_0 => "001010101100010101", xin_1 => "000101000100100110", pass => true),
  (xin_0 => "001101110011001100", xin_1 => "001001001011111111", pass => true),
  (xin_0 => "000111000000010000", xin_1 => "000101101100001001", pass => true),
  (xin_0 => "001001111100000111", xin_1 => "000010001001000111", pass => false),
  (xin_0 => "001011011000100101", xin_1 => "000010101110011111", pass => true),
  (xin_0 => "001000000101101110", xin_1 => "000110101101011000", pass => true),
  (xin_0 => "000101011100110010", xin_1 => "000100000000000011", pass => true),
  (xin_0 => "001001111010101001", xin_1 => "000100101000000001", pass => true),
  (xin_0 => "001001101010110100", xin_1 => "000010010110011010", pass => false),
  (xin_0 => "001000000001010001", xin_1 => "000111110110100011", pass => true),
  (xin_0 => "000100110101001000", xin_1 => "001001101011001111", pass => false),
  (xin_0 => "001111111111100101", xin_1 => "001000110111100110", pass => true),
  (xin_0 => "000111101011100111", xin_1 => "000011010011101100", pass => false),
  (xin_0 => "001011100001001001", xin_1 => "000101000110001001", pass => true),
  (xin_0 => "000111110010011010", xin_1 => "000010110110000001", pass => false),
  (xin_0 => "001000101000100110", xin_1 => "000010100011100110", pass => false),
  (xin_0 => "001001111000000001", xin_1 => "000011100101010110", pass => false),
  (xin_0 => "001100100010110000", xin_1 => "000111010001000011", pass => false),
  (xin_0 => "000111001011000000", xin_1 => "000011010001111010", pass => false),
  (xin_0 => "001001101111010101", xin_1 => "000111011000100010", pass => true),
  (xin_0 => "001000110001110010", xin_1 => "001011001111001111", pass => false),
  (xin_0 => "000111011110101011", xin_1 => "001000111111111100", pass => false),
  (xin_0 => "001001110110000011", xin_1 => "000011011100111110", pass => false),
  (xin_0 => "000101100011001001", xin_1 => "000110101100111111", pass => true),
  (xin_0 => "001011111101001011", xin_1 => "001000101101010111", pass => false),
  (xin_0 => "001000011011001100", xin_1 => "000001100010101111", pass => false),
  (xin_0 => "001001000101111101", xin_1 => "001000110111000101", pass => false),
  (xin_0 => "000111011001100011", xin_1 => "001001101010000111", pass => false),
  (xin_0 => "000111111110000011", xin_1 => "001000101011010101", pass => true),
  (xin_0 => "001001101011110000", xin_1 => "000111000000110100", pass => true),
  (xin_0 => "001100010111100011", xin_1 => "000111011010110101", pass => false),
  (xin_0 => "000111100001001101", xin_1 => "000010100101001100", pass => false),
  (xin_0 => "001001000011000010", xin_1 => "000001110010000001", pass => false),
  (xin_0 => "000101010011000100", xin_1 => "000100110101101011", pass => true),
  (xin_0 => "010000011010001101", xin_1 => "001001001110111010", pass => true),
  (xin_0 => "001001100000000101", xin_1 => "001010010101101010", pass => false),
  (xin_0 => "001011101010001010", xin_1 => "000111010100001100", pass => false),
  (xin_0 => "001000011110110001", xin_1 => "000101000001001011", pass => true),
  (xin_0 => "001011000101010111", xin_1 => "001001000011110010", pass => false),
  (xin_0 => "000100111000111001", xin_1 => "000110111110100100", pass => true),
  (xin_0 => "001000011010110101", xin_1 => "000110001000011101", pass => true),
  (xin_0 => "001001000111000100", xin_1 => "000011010010011001", pass => false),
  (xin_0 => "001000111011010000", xin_1 => "000101001101001010", pass => true),
  (xin_0 => "001101111000110110", xin_1 => "000110001111000000", pass => false),
  (xin_0 => "001000111101110011", xin_1 => "001011000111000011", pass => false),
  (xin_0 => "000101111101101101", xin_1 => "000100111100011111", pass => true),
  (xin_0 => "000111110110010100", xin_1 => "000011011100000110", pass => false),
  (xin_0 => "000111101111111000", xin_1 => "000110111110011011", pass => true),
  (xin_0 => "001000001101110101", xin_1 => "000010000100011101", pass => false),
  (xin_0 => "001010011101000011", xin_1 => "001011011001111111", pass => false),
  (xin_0 => "001100111100010101", xin_1 => "001000100000001100", pass => false),
  (xin_0 => "000111011100101101", xin_1 => "000011001011010100", pass => false),
  (xin_0 => "000110000001001001", xin_1 => "001001011111100001", pass => false),
  (xin_0 => "000100001111100111", xin_1 => "000010001110100000", pass => true),
  (xin_0 => "000111011011011100", xin_1 => "001010000011001110", pass => false),
  (xin_0 => "001011000011100010", xin_1 => "001010011100101111", pass => false),
  (xin_0 => "001101101011010010", xin_1 => "000100100101101011", pass => false),
  (xin_0 => "001110000101100110", xin_1 => "000110010001000110", pass => false),
  (xin_0 => "001100100000011100", xin_1 => "000111010011011010", pass => false),
  (xin_0 => "001111100101010010", xin_1 => "001001111011001000", pass => true),
  (xin_0 => "001011111010101010", xin_1 => "000100000000110110", pass => true),
  (xin_0 => "001110001011001011", xin_1 => "001000100001110000", pass => false),
  (xin_0 => "001001101100101011", xin_1 => "000110101100011111", pass => true),
  (xin_0 => "001011001001010001", xin_1 => "000110000000110001", pass => true),
  (xin_0 => "001011000101000110", xin_1 => "000101100101010011", pass => true),
  (xin_0 => "001010000001011100", xin_1 => "000111101101111001", pass => true),
  (xin_0 => "001011101010010010", xin_1 => "000111001100110001", pass => false),
  (xin_0 => "001000100111100111", xin_1 => "000100000010101011", pass => false),
  (xin_0 => "000101101110011011", xin_1 => "000111000100001110", pass => true),
  (xin_0 => "001101110001100100", xin_1 => "000101000000010101", pass => false),
  (xin_0 => "001101001000101000", xin_1 => "000110000101110111", pass => false),
  (xin_0 => "000110101100100110", xin_1 => "001000010010000011", pass => true),
  (xin_0 => "001011000010010111", xin_1 => "001000100010001110", pass => false),
  (xin_0 => "001100100100010101", xin_1 => "000001010011100101", pass => true),
  (xin_0 => "001010110010001011", xin_1 => "001011100001000001", pass => false),
  (xin_0 => "001100111000011100", xin_1 => "001000110101110111", pass => false),
  (xin_0 => "001100010100110000", xin_1 => "000011111001000110", pass => true),
  (xin_0 => "001001100000011001", xin_1 => "000010010010110010", pass => false),
  (xin_0 => "001100001101010101", xin_1 => "000111100000101011", pass => false),
  (xin_0 => "001100110010101011", xin_1 => "000111010111110011", pass => false),
  (xin_0 => "001011000100101110", xin_1 => "000111101110100001", pass => false),
  (xin_0 => "000111001101001101", xin_1 => "001010001100001111", pass => false),
  (xin_0 => "001011010110000001", xin_1 => "000010010100110100", pass => true),
  (xin_0 => "001000001010111110", xin_1 => "000110010000110101", pass => true),
  (xin_0 => "000100100100111101", xin_1 => "000010000000010110", pass => true),
  (xin_0 => "000111000011101011", xin_1 => "000011001100001100", pass => false),
  (xin_0 => "001001011110110101", xin_1 => "000101111110100011", pass => true),
  (xin_0 => "000100110011101001", xin_1 => "000110010100000010", pass => true),
  (xin_0 => "000110011000000101", xin_1 => "000100111101011010", pass => true),
  (xin_0 => "000101110110101000", xin_1 => "001010001100011001", pass => false),
  (xin_0 => "001011100101011111", xin_1 => "000111110100000011", pass => false),
  (xin_0 => "001001011001001000", xin_1 => "001010111000101000", pass => false),
  (xin_0 => "000111110111100000", xin_1 => "001010011000000011", pass => false),
  (xin_0 => "001101001101111010", xin_1 => "001001111001001000", pass => true),
  (xin_0 => "000111110001111100", xin_1 => "000010111010100011", pass => false),
  (xin_0 => "001010000011100110", xin_1 => "001010111100100101", pass => false),
  (xin_0 => "001011111101100010", xin_1 => "001001000011011010", pass => false),
  (xin_0 => "001101010011101010", xin_1 => "000101000100101101", pass => false),
  (xin_0 => "001000011101110010", xin_1 => "001010001111011100", pass => false),
  (xin_0 => "001001011101010100", xin_1 => "001100000100110001", pass => false),
  (xin_0 => "001001101010010001", xin_1 => "000100001000010010", pass => true),
  (xin_0 => "001011001011011001", xin_1 => "000010011011101001", pass => true),
  (xin_0 => "001001100101010110", xin_1 => "000101000110111011", pass => true),
  (xin_0 => "000111001110100010", xin_1 => "000010001010111010", pass => false),
  (xin_0 => "001000011110011101", xin_1 => "000100000110111100", pass => false),
  (xin_0 => "001010101100110001", xin_1 => "000101111001101000", pass => true),
  (xin_0 => "001011000001011011", xin_1 => "000010111011111111", pass => true),
  (xin_0 => "000010111000011000", xin_1 => "000100011001000000", pass => true),
  (xin_0 => "000101101111111100", xin_1 => "000101001010010011", pass => true),
  (xin_0 => "001010101011110110", xin_1 => "001000110100111111", pass => false),
  (xin_0 => "000111000000010111", xin_1 => "001000010011011010", pass => true),
  (xin_0 => "001010011001000110", xin_1 => "001010000100110010", pass => false),
  (xin_0 => "001101111100001101", xin_1 => "000100110111011000", pass => false),
  (xin_0 => "001100000010001111", xin_1 => "000100001000010011", pass => true),
  (xin_0 => "001001110001001110", xin_1 => "000001111000000011", pass => false),
  (xin_0 => "000110100110100001", xin_1 => "000010100011110010", pass => false),
  (xin_0 => "000110101010010011", xin_1 => "000001110101110110", pass => false),
  (xin_0 => "000100111110100111", xin_1 => "001001001010111000", pass => false),
  (xin_0 => "001100011110101001", xin_1 => "000110111110100010", pass => false),
  (xin_0 => "001011101100100101", xin_1 => "000011100001111000", pass => true),
  (xin_0 => "000011000011110100", xin_1 => "000010011110101110", pass => true),
  (xin_0 => "000111001101111010", xin_1 => "001010100111100110", pass => false),
  (xin_0 => "001101010001011001", xin_1 => "000001100100010000", pass => true),
  (xin_0 => "000110111010011011", xin_1 => "001010101010101011", pass => false),
  (xin_0 => "001001001000001101", xin_1 => "001011001110010111", pass => false),
  (xin_0 => "000111110001011100", xin_1 => "001000000011101110", pass => true),
  (xin_0 => "001101110011111001", xin_1 => "000110100100011111", pass => false),
  (xin_0 => "001101001010001011", xin_1 => "000101011011111111", pass => false),
  (xin_0 => "000010010101011001", xin_1 => "000011001000010101", pass => true),
  (xin_0 => "001010110110100110", xin_1 => "001010000000110110", pass => false),
  (xin_0 => "001000011010001111", xin_1 => "000010010111110001", pass => false),
  (xin_0 => "001110001010100101", xin_1 => "001010111000011110", pass => true),
  (xin_0 => "001000001110111111", xin_1 => "000111110010101001", pass => true),
  (xin_0 => "000111001110110111", xin_1 => "001010000000100001", pass => false),
  (xin_0 => "001101000010001100", xin_1 => "000111001100101000", pass => false),
  (xin_0 => "001010001011110101", xin_1 => "000110010111011001", pass => true),
  (xin_0 => "000110100111100000", xin_1 => "001001000101101011", pass => false),
  (xin_0 => "000110001011110010", xin_1 => "000001010100101101", pass => false),
  (xin_0 => "001011111100011001", xin_1 => "001000100011100000", pass => false),
  (xin_0 => "001001100110101101", xin_1 => "001010010011011101", pass => false),
  (xin_0 => "010000010000011101", xin_1 => "001010100011111100", pass => true),
  (xin_0 => "001000100101011001", xin_1 => "000010001010111011", pass => false),
  (xin_0 => "000100111010111001", xin_1 => "000011010111001001", pass => true),
  (xin_0 => "000110100011101110", xin_1 => "000100101100000010", pass => true),
  (xin_0 => "001001011100000111", xin_1 => "000111010001110000", pass => true),
  (xin_0 => "010001000110101111", xin_1 => "001010001011110011", pass => true),
  (xin_0 => "000110001011001110", xin_1 => "000111011110011010", pass => true),
  (xin_0 => "000101011111101001", xin_1 => "000101001110110010", pass => true),
  (xin_0 => "001000001011001001", xin_1 => "001010011001001110", pass => false),
  (xin_0 => "001010111011011011", xin_1 => "001010110011001100", pass => false),
  (xin_0 => "001000101011101001", xin_1 => "000010010110001000", pass => false),
  (xin_0 => "000110110101001010", xin_1 => "000010001010010001", pass => false),
  (xin_0 => "000100001010110010", xin_1 => "000000000000100101", pass => true),
  (xin_0 => "001011101101011111", xin_1 => "000000011101001101", pass => true),
  (xin_0 => "000101101100111000", xin_1 => "000101010100111000", pass => true),
  (xin_0 => "001011110011111110", xin_1 => "000111000000110011", pass => false),
  (xin_0 => "001111111101001000", xin_1 => "001010110001100010", pass => true),
  (xin_0 => "000101011111110111", xin_1 => "000011110111111011", pass => true),
  (xin_0 => "000110111111001010", xin_1 => "000111110110110100", pass => true),
  (xin_0 => "001001110010010001", xin_1 => "000100101010000100", pass => true),
  (xin_0 => "000111000110011011", xin_1 => "000111110100000110", pass => true),
  (xin_0 => "010000011110001001", xin_1 => "000010101101111100", pass => false),
  (xin_0 => "010000110011101000", xin_1 => "001010010100100010", pass => true),
  (xin_0 => "001010010000110111", xin_1 => "000101100110111010", pass => true),
  (xin_0 => "000110110011111111", xin_1 => "000111111110111101", pass => true),
  (xin_0 => "000111001001111000", xin_1 => "000010110101010111", pass => false),
  (xin_0 => "001011101101110000", xin_1 => "001000011010011010", pass => false),
  (xin_0 => "001001000011000110", xin_1 => "001011111011111110", pass => false),
  (xin_0 => "001111110011010111", xin_1 => "001010010001011011", pass => true),
  (xin_0 => "000111000001101100", xin_1 => "001011000111101001", pass => false),
  (xin_0 => "001101010001000000", xin_1 => "000111011001100011", pass => false),
  (xin_0 => "000101111110010100", xin_1 => "000101001001000100", pass => true),
  (xin_0 => "000111010100000101", xin_1 => "000001010011001111", pass => false),
  (xin_0 => "001000001100100110", xin_1 => "000010010111011101", pass => false),
  (xin_0 => "001100000011110001", xin_1 => "001000000101010010", pass => false),
  (xin_0 => "000110111100011111", xin_1 => "001001000111111010", pass => false),
  (xin_0 => "001011001011110110", xin_1 => "001010011110100000", pass => false),
  (xin_0 => "001011101011100110", xin_1 => "000101011101001010", pass => true),
  (xin_0 => "000101011111010111", xin_1 => "001001000001100001", pass => false),
  (xin_0 => "000110110000101010", xin_1 => "000111001000100111", pass => true),
  (xin_0 => "001010000100100011", xin_1 => "001100000011001000", pass => false),
  (xin_0 => "000110110011010000", xin_1 => "001000010011110100", pass => true),
  (xin_0 => "001011010111010111", xin_1 => "000010010010101111", pass => true),
  (xin_0 => "001011100100011100", xin_1 => "000010101011101101", pass => true),
  (xin_0 => "001011011011100101", xin_1 => "001001001001000011", pass => false),
  (xin_0 => "001101000010010100", xin_1 => "111111110111001110", pass => true),
  (xin_0 => "000110110111011110", xin_1 => "000110110011010101", pass => true),
  (xin_0 => "000111100110001100", xin_1 => "000101100110100100", pass => true),
  (xin_0 => "000101110111010000", xin_1 => "000111000000011011", pass => true),
  (xin_0 => "000111110100111111", xin_1 => "000010111011100001", pass => false),
  (xin_0 => "000110100011000011", xin_1 => "000010111100110100", pass => false),
  (xin_0 => "001010100111000100", xin_1 => "000011110000101010", pass => true),
  (xin_0 => "001100010000001000", xin_1 => "000001011100100111", pass => true),
  (xin_0 => "001001100000111001", xin_1 => "000010011000000100", pass => false),
  (xin_0 => "000111111110011100", xin_1 => "000001110100010000", pass => false),
  (xin_0 => "001000010101010100", xin_1 => "000010010110110100", pass => false),
  (xin_0 => "000110101000100110", xin_1 => "000101010111101101", pass => true),
  (xin_0 => "001011010111010010", xin_1 => "000111100100100010", pass => false),
  (xin_0 => "001011100110101111", xin_1 => "001000000101011010", pass => false),
  (xin_0 => "001010101111111010", xin_1 => "000011001110101100", pass => true),
  (xin_0 => "001001010111100111", xin_1 => "000111010000001110", pass => true),
  (xin_0 => "000100111010111100", xin_1 => "000100001010010101", pass => true),
  (xin_0 => "000011000110001000", xin_1 => "000011110100100001", pass => true),
  (xin_0 => "001001010011010010", xin_1 => "000010110101001000", pass => false),
  (xin_0 => "001010111010110010", xin_1 => "001001001001100000", pass => false),
  (xin_0 => "001101001110000110", xin_1 => "000111111110010010", pass => false),
  (xin_0 => "001011010011100101", xin_1 => "001000011000011000", pass => false),
  (xin_0 => "000111111010100101", xin_1 => "000011000111100111", pass => false),
  (xin_0 => "001101001100001011", xin_1 => "000101111000111110", pass => false),
  (xin_0 => "000011000011000001", xin_1 => "000011010000010100", pass => true),
  (xin_0 => "001000010111110011", xin_1 => "000111000110011101", pass => true),
  (xin_0 => "000100111100100000", xin_1 => "000110100001011111", pass => true),
  (xin_0 => "001001001110011101", xin_1 => "001010100111000001", pass => false),
  (xin_0 => "001110010111110011", xin_1 => "001001101011001101", pass => true),
  (xin_0 => "001000100100000010", xin_1 => "000010110011101100", pass => false),
  (xin_0 => "000111100001011000", xin_1 => "000010100001101010", pass => false),
  (xin_0 => "001010011100001100", xin_1 => "001000011110110000", pass => false),
  (xin_0 => "000110111010110100", xin_1 => "000011110000101101", pass => false),
  (xin_0 => "001010010110000100", xin_1 => "000010101110011101", pass => false),
  (xin_0 => "001000111110101000", xin_1 => "001010101100100101", pass => false),
  (xin_0 => "000101101001101111", xin_1 => "000100101110011010", pass => true),
  (xin_0 => "001011010111100000", xin_1 => "000100011011010001", pass => true),
  (xin_0 => "001011110101101001", xin_1 => "001001011000110010", pass => false),
  (xin_0 => "000110110110011100", xin_1 => "000010101011010011", pass => false),
  (xin_0 => "001001111100010011", xin_1 => "000010001101011111", pass => false),
  (xin_0 => "000011111011100010", xin_1 => "000111111011111100", pass => false),
  (xin_0 => "001000000010110001", xin_1 => "000110010010010110", pass => true),
  (xin_0 => "001010010010110100", xin_1 => "001001000100100001", pass => false),
  (xin_0 => "000000101111000100", xin_1 => "000101101100000111", pass => false),
  (xin_0 => "001011010101101011", xin_1 => "000101011110010101", pass => true),
  (xin_0 => "001100100011110101", xin_1 => "001010101001010111", pass => true),
  (xin_0 => "000101010110011100", xin_1 => "000101001010001000", pass => true),
  (xin_0 => "001010001110101001", xin_1 => "000011011000100000", pass => false),
  (xin_0 => "000101000011101011", xin_1 => "001000101011001000", pass => false),
  (xin_0 => "000110000001011000", xin_1 => "001000100011111011", pass => false),
  (xin_0 => "001000111000001010", xin_1 => "000010000010101111", pass => false),
  (xin_0 => "001000000110010011", xin_1 => "000010100000011000", pass => false),
  (xin_0 => "001100111011100100", xin_1 => "000111100001110010", pass => false),
  (xin_0 => "001010011100111111", xin_1 => "001010100000001011", pass => false),
  (xin_0 => "001011101111001000", xin_1 => "000011011111011101", pass => true),
  (xin_0 => "001000100011101001", xin_1 => "000001111111100100", pass => false),
  (xin_0 => "001011011111010000", xin_1 => "000001110000110111", pass => true),
  (xin_0 => "001000101110010111", xin_1 => "000110111010101110", pass => true),
  (xin_0 => "000100000001011011", xin_1 => "000100011111110110", pass => true),
  (xin_0 => "000111010100110110", xin_1 => "000011001001100100", pass => false),
  (xin_0 => "000111100101001000", xin_1 => "000011011101010110", pass => false),
  (xin_0 => "001100101100001011", xin_1 => "000100001110110011", pass => true),
  (xin_0 => "001011000010111100", xin_1 => "000111010110001100", pass => false),
  (xin_0 => "001011001101000010", xin_1 => "000111001011010101", pass => false),
  (xin_0 => "001001110101010011", xin_1 => "001011000111010001", pass => false),
  (xin_0 => "001010011101111000", xin_1 => "001010101010100110", pass => false),
  (xin_0 => "001100010101000011", xin_1 => "000111100101010110", pass => false),
  (xin_0 => "000101111111100000", xin_1 => "001000111010010110", pass => false),
  (xin_0 => "001000101100110011", xin_1 => "000011010110001000", pass => false),
  (xin_0 => "001011101000010011", xin_1 => "001000010110111111", pass => false),
  (xin_0 => "000101111100110001", xin_1 => "001001011001011100", pass => false),
  (xin_0 => "000110011000110100", xin_1 => "001001011011100111", pass => false),
  (xin_0 => "000011100001111000", xin_1 => "000010101011010101", pass => true),
  (xin_0 => "001100010010000100", xin_1 => "001000001001111101", pass => false),
  (xin_0 => "001011110111100011", xin_1 => "000010110100110011", pass => true),
  (xin_0 => "000111010010110110", xin_1 => "001001110000010001", pass => false),
  (xin_0 => "001011010001100101", xin_1 => "000100010010001111", pass => true),
  (xin_0 => "000100000110101110", xin_1 => "001000010001010100", pass => false),
  (xin_0 => "001010110111011011", xin_1 => "001000110001000001", pass => false),
  (xin_0 => "000110001001100000", xin_1 => "000101100010100001", pass => true),
  (xin_0 => "001001010011011011", xin_1 => "001011011101101000", pass => false),
  (xin_0 => "001001010011111000", xin_1 => "000010011100111100", pass => false),
  (xin_0 => "001100010110011101", xin_1 => "000100100000010110", pass => true),
  (xin_0 => "001100000100001001", xin_1 => "000010000010100010", pass => true),
  (xin_0 => "001010000101001100", xin_1 => "000011110010000100", pass => true),
  (xin_0 => "001011010010111111", xin_1 => "001000011110101010", pass => false),
  (xin_0 => "001100001100111101", xin_1 => "000110110000010001", pass => false),
  (xin_0 => "001000110011001111", xin_1 => "000011111101011101", pass => false),
  (xin_0 => "001100100010000101", xin_1 => "000111100100011001", pass => false),
  (xin_0 => "001110111001101111", xin_1 => "000101111010000111", pass => false),
  (xin_0 => "000101000001011011", xin_1 => "000101011100011000", pass => true),
  (xin_0 => "000111101100001100", xin_1 => "001010101000011010", pass => false),
  (xin_0 => "001000100011110110", xin_1 => "000001111011010100", pass => false),
  (xin_0 => "001000000011101110", xin_1 => "001001110000110000", pass => false),
  (xin_0 => "001010010110110000", xin_1 => "001001011000000100", pass => false),
  (xin_0 => "001001110111010010", xin_1 => "001010111010001001", pass => false),
  (xin_0 => "001001011001001010", xin_1 => "000011010011000011", pass => false),
  (xin_0 => "000110111000100100", xin_1 => "000001001100111100", pass => false),
  (xin_0 => "001000101111000010", xin_1 => "000111000010011011", pass => true),
  (xin_0 => "001011110110001100", xin_1 => "001000101100010111", pass => false),
  (xin_0 => "001100110110111100", xin_1 => "001000010010001110", pass => false),
  (xin_0 => "000100110000111000", xin_1 => "000010100000101100", pass => true),
  (xin_0 => "001010100011000110", xin_1 => "001000110101010011", pass => false),
  (xin_0 => "001101001001010111", xin_1 => "000110110111100010", pass => false),
  (xin_0 => "001100000111001001", xin_1 => "000010111001000011", pass => true),
  (xin_0 => "001000101110101011", xin_1 => "000010100001011011", pass => false),
  (xin_0 => "000110011011010000", xin_1 => "000111000001000110", pass => true),
  (xin_0 => "000011001001110110", xin_1 => "000111011101000011", pass => false),
  (xin_0 => "000100110010100011", xin_1 => "000011110111110001", pass => true),
  (xin_0 => "000111000001111000", xin_1 => "001001110100101110", pass => false),
  (xin_0 => "001100110000011111", xin_1 => "000010111100000000", pass => true),
  (xin_0 => "001001011100101100", xin_1 => "000100101100110111", pass => true),
  (xin_0 => "000101111111110001", xin_1 => "000001111000111101", pass => false),
  (xin_0 => "001011100111000010", xin_1 => "000111110100101010", pass => false),
  (xin_0 => "001000010000101010", xin_1 => "000100010110001011", pass => false),
  (xin_0 => "001011101011011100", xin_1 => "000011110101000100", pass => true),
  (xin_0 => "001010000100111001", xin_1 => "001011011100101110", pass => false),
  (xin_0 => "001000010101111100", xin_1 => "000101001101100110", pass => true),
  (xin_0 => "000110111001011100", xin_1 => "000011010111001110", pass => false),
  (xin_0 => "001101101001011001", xin_1 => "000110001010111011", pass => false),
  (xin_0 => "000101000100010110", xin_1 => "000110101010111110", pass => true),
  (xin_0 => "001100001100100010", xin_1 => "000010100001110010", pass => true),
  (xin_0 => "000100110101110101", xin_1 => "000110000000000010", pass => true),
  (xin_0 => "000111000101110110", xin_1 => "001011010110010011", pass => false),
  (xin_0 => "001001110111100101", xin_1 => "000100011001101110", pass => true),
  (xin_0 => "000100101010111100", xin_1 => "000101010100110110", pass => true),
  (xin_0 => "000111100100011101", xin_1 => "000010011100010010", pass => false),
  (xin_0 => "000010110101110101", xin_1 => "000110110100000010", pass => false),
  (xin_0 => "001100010110011010", xin_1 => "001000110111011101", pass => false),
  (xin_0 => "000111111011000110", xin_1 => "001010000110101010", pass => false),
  (xin_0 => "001110010011101001", xin_1 => "000101000101010000", pass => false),
  (xin_0 => "001011100110100111", xin_1 => "001001101101101001", pass => false),
  (xin_0 => "001000000001010101", xin_1 => "000010110100110010", pass => false),
  (xin_0 => "001101000000011010", xin_1 => "000111100010010011", pass => false),
  (xin_0 => "001011011101000111", xin_1 => "001000100011010110", pass => false),
  (xin_0 => "001001011101010110", xin_1 => "000010110111011111", pass => false),
  (xin_0 => "000111010100110110", xin_1 => "000010110101011101", pass => false),
  (xin_0 => "000110001001001000", xin_1 => "000001010110101101", pass => false),
  (xin_0 => "001000111001110000", xin_1 => "000010100010011000", pass => false),
  (xin_0 => "001101001110000001", xin_1 => "000110000011010100", pass => false),
  (xin_0 => "000111100110100011", xin_1 => "000011101001000100", pass => false),
  (xin_0 => "001000001001000001", xin_1 => "000010010010000111", pass => false),
  (xin_0 => "000011100100010100", xin_1 => "000011010000011010", pass => true),
  (xin_0 => "001000000101110000", xin_1 => "000011101110010111", pass => false),
  (xin_0 => "000101101011010110", xin_1 => "001000000011010000", pass => false),
  (xin_0 => "001011110100101110", xin_1 => "000010111000011111", pass => true),
  (xin_0 => "001001000100000010", xin_1 => "000001001111110011", pass => false),
  (xin_0 => "000101001001000011", xin_1 => "000101111101011100", pass => true),
  (xin_0 => "001100011111000011", xin_1 => "001001011000001111", pass => false),
  (xin_0 => "001011101111000000", xin_1 => "000100101000111101", pass => true),
  (xin_0 => "001100001011101111", xin_1 => "000111100001110010", pass => false),
  (xin_0 => "000101100000111110", xin_1 => "001000101100111011", pass => false),
  (xin_0 => "001100111100010110", xin_1 => "000100010001000110", pass => true),
  (xin_0 => "001001110000001011", xin_1 => "000101100100001110", pass => true),
  (xin_0 => "001010100001111010", xin_1 => "000011101010101111", pass => true),
  (xin_0 => "000100000101110001", xin_1 => "001001100000001110", pass => false),
  (xin_0 => "001010000100010010", xin_1 => "001100110001101100", pass => false),
  (xin_0 => "000101011100000011", xin_1 => "001001000001001100", pass => false),
  (xin_0 => "000100000011100011", xin_1 => "000101101100001111", pass => true),
  (xin_0 => "001100010100101011", xin_1 => "001000001101110001", pass => false),
  (xin_0 => "001011100011100100", xin_1 => "000100000010101100", pass => true),
  (xin_0 => "001010010100010011", xin_1 => "001100011001010011", pass => false),
  (xin_0 => "000110110001011011", xin_1 => "000101010000000010", pass => true),
  (xin_0 => "000111110101001110", xin_1 => "000110100010110101", pass => true),
  (xin_0 => "001000001111000001", xin_1 => "000001000101111101", pass => false),
  (xin_0 => "000101000111101001", xin_1 => "000101110010000111", pass => true),
  (xin_0 => "001101001100011001", xin_1 => "000110011011100000", pass => false),
  (xin_0 => "000111110000000101", xin_1 => "000111101000100111", pass => true),
  (xin_0 => "001100011010100010", xin_1 => "001000101100011111", pass => false),
  (xin_0 => "000101100010100010", xin_1 => "000101111011100010", pass => true),
  (xin_0 => "000101111111000110", xin_1 => "000011001001110110", pass => false),
  (xin_0 => "000111001100101011", xin_1 => "000101110101011001", pass => true),
  (xin_0 => "001100110000011000", xin_1 => "000110110110111100", pass => false),
  (xin_0 => "001010000011001010", xin_1 => "001001001110100001", pass => false),
  (xin_0 => "000110100100001100", xin_1 => "001000110101100000", pass => false),
  (xin_0 => "001010000111110110", xin_1 => "000010111000110000", pass => false),
  (xin_0 => "001000011100000111", xin_1 => "000001110011111000", pass => false),
  (xin_0 => "000110100010000011", xin_1 => "001001001001000011", pass => false),
  (xin_0 => "001000000110000011", xin_1 => "000111110111001110", pass => true),
  (xin_0 => "000101111100011000", xin_1 => "000010011101101110", pass => false),
  (xin_0 => "000100011101000010", xin_1 => "000011001000110100", pass => true),
  (xin_0 => "001011010101000111", xin_1 => "000100101010100000", pass => true),
  (xin_0 => "000110000100100011", xin_1 => "000100101100000000", pass => true),
  (xin_0 => "000100011010011001", xin_1 => "001000001000110110", pass => false),
  (xin_0 => "001101101101100011", xin_1 => "001010111000111110", pass => true),
  (xin_0 => "001001101101010000", xin_1 => "001100000010110001", pass => false),
  (xin_0 => "000100100001110010", xin_1 => "000011001010000001", pass => true),
  (xin_0 => "000101010001011100", xin_1 => "000101011001100000", pass => true),
  (xin_0 => "001000000110000111", xin_1 => "000111000000000110", pass => true),
  (xin_0 => "001011011011110010", xin_1 => "000010110110101100", pass => true),
  (xin_0 => "001001001111011001", xin_1 => "000011000010001110", pass => false),
  (xin_0 => "000111011000010011", xin_1 => "000110001110100101", pass => true),
  (xin_0 => "000111010001111110", xin_1 => "000110110110101100", pass => true),
  (xin_0 => "000110000001011101", xin_1 => "000011111000101000", pass => true),
  (xin_0 => "000101101001001101", xin_1 => "001001000000100101", pass => false),
  (xin_0 => "001011010111100001", xin_1 => "001000001101100101", pass => false),
  (xin_0 => "001100111111000001", xin_1 => "000101000101011000", pass => false),
  (xin_0 => "000100010001010010", xin_1 => "000010101101100000", pass => true),
  (xin_0 => "000110101110110100", xin_1 => "000010010010000111", pass => false),
  (xin_0 => "000110000100011010", xin_1 => "000011011000010000", pass => false),
  (xin_0 => "000011001110000011", xin_1 => "000111010001100111", pass => false),
  (xin_0 => "001001001001010001", xin_1 => "001011001001110111", pass => false),
  (xin_0 => "000101101000011100", xin_1 => "000100101011110000", pass => true),
  (xin_0 => "000111111001111000", xin_1 => "000001000011001111", pass => false),
  (xin_0 => "001100010001011110", xin_1 => "001000101110110101", pass => false),
  (xin_0 => "000110100011100000", xin_1 => "000011101110111101", pass => false),
  (xin_0 => "000111000110000001", xin_1 => "000010001000000001", pass => false),
  (xin_0 => "001000001001001100", xin_1 => "000010111111111100", pass => false),
  (xin_0 => "000011010100001110", xin_1 => "000101101111100000", pass => true),
  (xin_0 => "001010110100110111", xin_1 => "000011011001010001", pass => true),
  (xin_0 => "000100010010001110", xin_1 => "000101000010101011", pass => true),
  (xin_0 => "000111000001101001", xin_1 => "000111010100000010", pass => true),
  (xin_0 => "000111110010110111", xin_1 => "000010101110110010", pass => false),
  (xin_0 => "000111000110100011", xin_1 => "000011000100100100", pass => false),
  (xin_0 => "001000101010000110", xin_1 => "000010010000011001", pass => false),
  (xin_0 => "001010010111111111", xin_1 => "000110110100001110", pass => true),
  (xin_0 => "001010111110111111", xin_1 => "000111111100010101", pass => false),
  (xin_0 => "001011000011010101", xin_1 => "001000010111110111", pass => false),
  (xin_0 => "000100010010001000", xin_1 => "000100110110110101", pass => true),
  (xin_0 => "000111010111001000", xin_1 => "001001010110011010", pass => false),
  (xin_0 => "001000110110001001", xin_1 => "000010000111100100", pass => false),
  (xin_0 => "001010010011011110", xin_1 => "000111000101010000", pass => true),
  (xin_0 => "010000111011110100", xin_1 => "001010101100111011", pass => true),
  (xin_0 => "001100011010011100", xin_1 => "000110110011011111", pass => false),
  (xin_0 => "000100011101101110", xin_1 => "000111011001100101", pass => false),
  (xin_0 => "000110011110110010", xin_1 => "000010101010000001", pass => false),
  (xin_0 => "001001001001101000", xin_1 => "000011111010101000", pass => false),
  (xin_0 => "000011100010000011", xin_1 => "000011001011101111", pass => true),
  (xin_0 => "001100110010100011", xin_1 => "000001101111010111", pass => true),
  (xin_0 => "001010100111101111", xin_1 => "000101001011111100", pass => true),
  (xin_0 => "000110111001001110", xin_1 => "000110011101010101", pass => true),
  (xin_0 => "001000011101001000", xin_1 => "000010001111000010", pass => false),
  (xin_0 => "000011111010111011", xin_1 => "000111010101111001", pass => false),
  (xin_0 => "000110100110001101", xin_1 => "000100001101010000", pass => true),
  (xin_0 => "000110110000011000", xin_1 => "001000101000111101", pass => false),
  (xin_0 => "001111001110001010", xin_1 => "001001110000001000", pass => true),
  (xin_0 => "001011100000110011", xin_1 => "000011001011010100", pass => true),
  (xin_0 => "000101010001111101", xin_1 => "000100000101101001", pass => true),
  (xin_0 => "001001000110110001", xin_1 => "000010001110111110", pass => false),
  (xin_0 => "001001000101000000", xin_1 => "000110001010101100", pass => true),
  (xin_0 => "001010000110010110", xin_1 => "000111100000111100", pass => true),
  (xin_0 => "000100100010101001", xin_1 => "000011111110100100", pass => true),
  (xin_0 => "001001110001000100", xin_1 => "000111010001011000", pass => true),
  (xin_0 => "000110010100010000", xin_1 => "000100011000011101", pass => true),
  (xin_0 => "000111110111011010", xin_1 => "000010000000011010", pass => false),
  (xin_0 => "000110011000010000", xin_1 => "000001011010000110", pass => false),
  (xin_0 => "001011011000010101", xin_1 => "001010110010011000", pass => false),
  (xin_0 => "001000100000110111", xin_1 => "000100001100011110", pass => false),
  (xin_0 => "000110011111000000", xin_1 => "000100011011110001", pass => true),
  (xin_0 => "000110101000111111", xin_1 => "000010100011100010", pass => false),
  (xin_0 => "001011110000101101", xin_1 => "001001000001110010", pass => false),
  (xin_0 => "000011011111110011", xin_1 => "000100110110001110", pass => true),
  (xin_0 => "001000101100001101", xin_1 => "001100010101111111", pass => false),
  (xin_0 => "001000001110110110", xin_1 => "000111110000110011", pass => true),
  (xin_0 => "001000101100111010", xin_1 => "000010001100100000", pass => false),
  (xin_0 => "001011000000111100", xin_1 => "001000100111100111", pass => false),
  (xin_0 => "000100000010101011", xin_1 => "001000000110000011", pass => false),
  (xin_0 => "001010010111000100", xin_1 => "001001011011001110", pass => false),
  (xin_0 => "001010001001111100", xin_1 => "000011001011011010", pass => false),
  (xin_0 => "001011010101110001", xin_1 => "000100001011101110", pass => true),
  (xin_0 => "000111001010000101", xin_1 => "000011001111000110", pass => false),
  (xin_0 => "000101100000000000", xin_1 => "001001111101010011", pass => false),
  (xin_0 => "001001010111100001", xin_1 => "001000110010111110", pass => false),
  (xin_0 => "000100101000100010", xin_1 => "000110111010111000", pass => true),
  (xin_0 => "000111010001010001", xin_1 => "000010010111011001", pass => false),
  (xin_0 => "001010000000101100", xin_1 => "001000001001100111", pass => false),
  (xin_0 => "000110101001110010", xin_1 => "001001111111101100", pass => false),
  (xin_0 => "001000100010000111", xin_1 => "000010000000101010", pass => false),
  (xin_0 => "000111110100100101", xin_1 => "001001100101001000", pass => false),
  (xin_0 => "000110010010101101", xin_1 => "000100011110001001", pass => true),
  (xin_0 => "000100100101000111", xin_1 => "000011010010100011", pass => true),
  (xin_0 => "001110011101000010", xin_1 => "000110000011100101", pass => false),
  (xin_0 => "001010010101001001", xin_1 => "000101000100100000", pass => true),
  (xin_0 => "000111100010000001", xin_1 => "001001111100110011", pass => false),
  (xin_0 => "000111110111101110", xin_1 => "000010111100101111", pass => false),
  (xin_0 => "000100100100111101", xin_1 => "000101011000110001", pass => true),
  (xin_0 => "001001101110001010", xin_1 => "000011000001001000", pass => false),
  (xin_0 => "000111101101010101", xin_1 => "000100000010001011", pass => false),
  (xin_0 => "000100100010000101", xin_1 => "000000111111010001", pass => true),
  (xin_0 => "000110110100100011", xin_1 => "000010110000101000", pass => false),
  (xin_0 => "001011011001100110", xin_1 => "001001111011000100", pass => false),
  (xin_0 => "001001110100111001", xin_1 => "000010010100010000", pass => false),
  (xin_0 => "001001100100101000", xin_1 => "000100110111000011", pass => true),
  (xin_0 => "001010110101101110", xin_1 => "001000011111010110", pass => false),
  (xin_0 => "000111111100001000", xin_1 => "000001101101100001", pass => false),
  (xin_0 => "000110011100001001", xin_1 => "001001100010001001", pass => false),
  (xin_0 => "000100000001000111", xin_1 => "000011101010001110", pass => true),
  (xin_0 => "000101110111111000", xin_1 => "001000001111111110", pass => false),
  (xin_0 => "001010101100001001", xin_1 => "001001101011011001", pass => false),
  (xin_0 => "001100100000011001", xin_1 => "000001111110111001", pass => true),
  (xin_0 => "000110101100100111", xin_1 => "000010110000000001", pass => false),
  (xin_0 => "000101001001101001", xin_1 => "000111101000100100", pass => false),
  (xin_0 => "001000010001100010", xin_1 => "000011010001000111", pass => false),
  (xin_0 => "000110001100011010", xin_1 => "000110001110101001", pass => true),
  (xin_0 => "000110110010011011", xin_1 => "000111101001101010", pass => true),
  (xin_0 => "001011000000100000", xin_1 => "001000111000001001", pass => false),
  (xin_0 => "001001011101011001", xin_1 => "000101001011100000", pass => true),
  (xin_0 => "001001111100010001", xin_1 => "000001111000101011", pass => false),
  (xin_0 => "000110001000011100", xin_1 => "001001011010101111", pass => false),
  (xin_0 => "001110000110011011", xin_1 => "000111000011011100", pass => false),
  (xin_0 => "001010000001100100", xin_1 => "000110000100100110", pass => true),
  (xin_0 => "001001001101101011", xin_1 => "000010111011001000", pass => false),
  (xin_0 => "000111111101101101", xin_1 => "000110011010101001", pass => true),
  (xin_0 => "001011101101101011", xin_1 => "000010010010000001", pass => true),
  (xin_0 => "000100100011000100", xin_1 => "000010011111110001", pass => true),
  (xin_0 => "000111100010111010", xin_1 => "000001100101010101", pass => false),
  (xin_0 => "000110011100100000", xin_1 => "001000100000101100", pass => false),
  (xin_0 => "001001101011011100", xin_1 => "000111101001001110", pass => true),
  (xin_0 => "001010101110110110", xin_1 => "000001110001100100", pass => false),
  (xin_0 => "000011110001101000", xin_1 => "000001110010111101", pass => true),
  (xin_0 => "000101110001001001", xin_1 => "000111011111111111", pass => true),
  (xin_0 => "001100000011010101", xin_1 => "001000001100010100", pass => false),
  (xin_0 => "001000110110101110", xin_1 => "000001001011010100", pass => false),
  (xin_0 => "000110000011100010", xin_1 => "000010100000010001", pass => false),
  (xin_0 => "000111001101111100", xin_1 => "000011010010110101", pass => false),
  (xin_0 => "001001101011110111", xin_1 => "000010010000101111", pass => false),
  (xin_0 => "001010101011111011", xin_1 => "000111101100101110", pass => false),
  (xin_0 => "001010011000111101", xin_1 => "000100010111000101", pass => true),
  (xin_0 => "000110000000000001", xin_1 => "000101010011010100", pass => true),
  (xin_0 => "001100001011111010", xin_1 => "000011111011100011", pass => true),
  (xin_0 => "001001010110111100", xin_1 => "000011110010111011", pass => false),
  (xin_0 => "000111011010111000", xin_1 => "000101001001001000", pass => true),
  (xin_0 => "001010000010011000", xin_1 => "000010000000011001", pass => false),
  (xin_0 => "001000101011101111", xin_1 => "001010110110011100", pass => false),
  (xin_0 => "000100100101111010", xin_1 => "000111000101100000", pass => true),
  (xin_0 => "001001001110100111", xin_1 => "000001011111001011", pass => false),
  (xin_0 => "001100011111111111", xin_1 => "000111110111110100", pass => false),
  (xin_0 => "001000110010010111", xin_1 => "000101100110000000", pass => true),
  (xin_0 => "001001000111101110", xin_1 => "000010001110001101", pass => false),
  (xin_0 => "000010000100110101", xin_1 => "000110001100100111", pass => false),
  (xin_0 => "001100011111000001", xin_1 => "000001011011101110", pass => true),
  (xin_0 => "001100010110001100", xin_1 => "000111011101110001", pass => false),
  (xin_0 => "000110110100111100", xin_1 => "000010111001100010", pass => false),
  (xin_0 => "000100011111111011", xin_1 => "000111110000010110", pass => false),
  (xin_0 => "001000000000111011", xin_1 => "000011000110110101", pass => false),
  (xin_0 => "001000011010001101", xin_1 => "000011001100011100", pass => false),
  (xin_0 => "001000110000010011", xin_1 => "001001000011101010", pass => false),
  (xin_0 => "001010111001100100", xin_1 => "001011000000011010", pass => false),
  (xin_0 => "000110110110101010", xin_1 => "000011010001010101", pass => false),
  (xin_0 => "000110010101111101", xin_1 => "000001011111001101", pass => false),
  (xin_0 => "001101001000100100", xin_1 => "000001100101111011", pass => true),
  (xin_0 => "001100001111110010", xin_1 => "000110101011010111", pass => false),
  (xin_0 => "001010100011001000", xin_1 => "001001000001110101", pass => false),
  (xin_0 => "001100111100000000", xin_1 => "001000111001001111", pass => false),
  (xin_0 => "001011000110110100", xin_1 => "000011001010100111", pass => true),
  (xin_0 => "000111011101010010", xin_1 => "001000110000001100", pass => true),
  (xin_0 => "001001100101010111", xin_1 => "001010001111101111", pass => false),
  (xin_0 => "001000111100011101", xin_1 => "000111110010010110", pass => true),
  (xin_0 => "000110101000101010", xin_1 => "000010000010110100", pass => false),
  (xin_0 => "001101111010000111", xin_1 => "000110010010110010", pass => false),
  (xin_0 => "000101001111011001", xin_1 => "000010111110011010", pass => true),
  (xin_0 => "001010011110101110", xin_1 => "001001110100111010", pass => false),
  (xin_0 => "000101100011100100", xin_1 => "001000000000100000", pass => false),
  (xin_0 => "001010001001110010", xin_1 => "000110101010000100", pass => true),
  (xin_0 => "000101101010001010", xin_1 => "001001110000100000", pass => false),
  (xin_0 => "000110000111000001", xin_1 => "000011000011111010", pass => false),
  (xin_0 => "001010010001110111", xin_1 => "000101110000000000", pass => true),
  (xin_0 => "000101001101101011", xin_1 => "000011000111000010", pass => true),
  (xin_0 => "001011010010010000", xin_1 => "000101100000011111", pass => true),
  (xin_0 => "001000110010110111", xin_1 => "000011000000101001", pass => false),
  (xin_0 => "001000111101001001", xin_1 => "000110000111011100", pass => true),
  (xin_0 => "001010001011100111", xin_1 => "000110011000111100", pass => true),
  (xin_0 => "000101011101000010", xin_1 => "000011110101111010", pass => true),
  (xin_0 => "001010011100000011", xin_1 => "000100101111001001", pass => true),
  (xin_0 => "001001001010011110", xin_1 => "000010001111010010", pass => false),
  (xin_0 => "001001111001010000", xin_1 => "000110110111111101", pass => true),
  (xin_0 => "001010100011010111", xin_1 => "000010111101101010", pass => true),
  (xin_0 => "001011111000010011", xin_1 => "000100111001100111", pass => true),
  (xin_0 => "000011110011111110", xin_1 => "001001010011111111", pass => false),
  (xin_0 => "000110011110111001", xin_1 => "000101011101001011", pass => true),
  (xin_0 => "000100110010011000", xin_1 => "000110100000011100", pass => true),
  (xin_0 => "001100001001100000", xin_1 => "000110111111110101", pass => false),
  (xin_0 => "001001110000000000", xin_1 => "000101100111010000", pass => true),
  (xin_0 => "001100110011000110", xin_1 => "001000101111000000", pass => false),
  (xin_0 => "001101011010111111", xin_1 => "000101001101010001", pass => false),
  (xin_0 => "000111011010100100", xin_1 => "000010011000000011", pass => false),
  (xin_0 => "000101001001100101", xin_1 => "000100101101101000", pass => true),
  (xin_0 => "001101001001111101", xin_1 => "000110111011000101", pass => false),
  (xin_0 => "001011111100001110", xin_1 => "001010001010000111", pass => false),
  (xin_0 => "000010110101010111", xin_1 => "000001110011110011", pass => true),
  (xin_0 => "000010111101100101", xin_1 => "000110010100110000", pass => false),
  (xin_0 => "001000000111001001", xin_1 => "001000010110101111", pass => true),
  (xin_0 => "001001100001000101", xin_1 => "000010010110101011", pass => false),
  (xin_0 => "000110110000110010", xin_1 => "000011010111000010", pass => false),
  (xin_0 => "001001001111010000", xin_1 => "001000001000110110", pass => true),
  (xin_0 => "001110000111110110", xin_1 => "001001010010000110", pass => true),
  (xin_0 => "001001000001011011", xin_1 => "000110011110110100", pass => true),
  (xin_0 => "001011000011100100", xin_1 => "000100010100111000", pass => true),
  (xin_0 => "001100110011011100", xin_1 => "001010110011111000", pass => true),
  (xin_0 => "001100011010101001", xin_1 => "000111001000100001", pass => false),
  (xin_0 => "001101001011111111", xin_1 => "000011000000010000", pass => true),
  (xin_0 => "001000111110111111", xin_1 => "000110010011100101", pass => true),
  (xin_0 => "000101110111011101", xin_1 => "000110010111011100", pass => true),
  (xin_0 => "000101110101000010", xin_1 => "000010101010010110", pass => false),
  (xin_0 => "000110011010100001", xin_1 => "000110111011101110", pass => true),
  (xin_0 => "000111111111000010", xin_1 => "000110110001100111", pass => true),
  (xin_0 => "000111101011111101", xin_1 => "000011110101000011", pass => false),
  (xin_0 => "001110111010001000", xin_1 => "001001100111101110", pass => true),
  (xin_0 => "001000111110101101", xin_1 => "000110001100111011", pass => true),
  (xin_0 => "010000000101111010", xin_1 => "001001111100111111", pass => true),
  (xin_0 => "001010011110000110", xin_1 => "000111000101100100", pass => true),
  (xin_0 => "001000001011100001", xin_1 => "001010011000011001", pass => false),
  (xin_0 => "001000110100011101", xin_1 => "001011001111010010", pass => false),
  (xin_0 => "001010100111101011", xin_1 => "000101101001100111", pass => true),
  (xin_0 => "000101100101111001", xin_1 => "000101010111001010", pass => true),
  (xin_0 => "000100100101011111", xin_1 => "000010101100100111", pass => true),
  (xin_0 => "001000110101011000", xin_1 => "000111001100110100", pass => true),
  (xin_0 => "001011111001000011", xin_1 => "000111111010100000", pass => false),
  (xin_0 => "000110101010010001", xin_1 => "000001111000100111", pass => false),
  (xin_0 => "000101101000000101", xin_1 => "000100100100011101", pass => true),
  (xin_0 => "000110100111000111", xin_1 => "000001101010100110", pass => false),
  (xin_0 => "001000110110000101", xin_1 => "000010001110100110", pass => false),
  (xin_0 => "000100100110000000", xin_1 => "000010110000101111", pass => true),
  (xin_0 => "001010001110011110", xin_1 => "001010110010001111", pass => false),
  (xin_0 => "001010000011100010", xin_1 => "000010001000010111", pass => false),
  (xin_0 => "001001000010111100", xin_1 => "000001101010011101", pass => false),
  (xin_0 => "001000101110110010", xin_1 => "000110001110100110", pass => true),
  (xin_0 => "001011010010000100", xin_1 => "001000000011010111", pass => false),
  (xin_0 => "001010111100101110", xin_1 => "000100101100000011", pass => true),
  (xin_0 => "001011100100100111", xin_1 => "001001001011010100", pass => false),
  (xin_0 => "001001000000111001", xin_1 => "000011010001010001", pass => false),
  (xin_0 => "001000000000010110", xin_1 => "001000000101100011", pass => true),
  (xin_0 => "001011100111111001", xin_1 => "000111001000111011", pass => false),
  (xin_0 => "001000100111111001", xin_1 => "000001101011011000", pass => false),
  (xin_0 => "001110011001010000", xin_1 => "000101000110111000", pass => false),
  (xin_0 => "000111001011001000", xin_1 => "000001111001010010", pass => false),
  (xin_0 => "001010101110001101", xin_1 => "000111101101100011", pass => false),
  (xin_0 => "001010110001010011", xin_1 => "000110000010010101", pass => true),
  (xin_0 => "000100001000001101", xin_1 => "000010011010000100", pass => true),
  (xin_0 => "001010001010111110", xin_1 => "001001100011101101", pass => false),
  (xin_0 => "000101000100111011", xin_1 => "000111110111100110", pass => false),
  (xin_0 => "000100101101101110", xin_1 => "001000001110010101", pass => false),
  (xin_0 => "000110011101001001", xin_1 => "000110000010101001", pass => true),
  (xin_0 => "001011101101000111", xin_1 => "000110001000110010", pass => true),
  (xin_0 => "000100111001011011", xin_1 => "000111101010111110", pass => false),
  (xin_0 => "000101101010011011", xin_1 => "000110010101001000", pass => true),
  (xin_0 => "000010101111100101", xin_1 => "000100110010000000", pass => true),
  (xin_0 => "001011010100110101", xin_1 => "000111111000101110", pass => false),
  (xin_0 => "000111001100011111", xin_1 => "000001010111110011", pass => false),
  (xin_0 => "000101010101100011", xin_1 => "000100001000100000", pass => true),
  (xin_0 => "000111000101100101", xin_1 => "000011110110111000", pass => false),
  (xin_0 => "000111011010001111", xin_1 => "001001111011010100", pass => false),
  (xin_0 => "000101010110001110", xin_1 => "000100101101110010", pass => true),
  (xin_0 => "001001011010101110", xin_1 => "000001111101010001", pass => false),
  (xin_0 => "001100000110011001", xin_1 => "001000101100011110", pass => false),
  (xin_0 => "001100000100101000", xin_1 => "001000010011100000", pass => false),
  (xin_0 => "000110001101011101", xin_1 => "000111100101000101", pass => true),
  (xin_0 => "000111110000110000", xin_1 => "001000011100000000", pass => true),
  (xin_0 => "001010011111111111", xin_1 => "001100110001011100", pass => false),
  (xin_0 => "000111101000111100", xin_1 => "000110000000001111", pass => true),
  (xin_0 => "001010110111100101", xin_1 => "001001110111010011", pass => false),
  (xin_0 => "001111110100001101", xin_1 => "001001101100001000", pass => true),
  (xin_0 => "001111000111010010", xin_1 => "001001101111100011", pass => true),
  (xin_0 => "000100001100001010", xin_1 => "000011010011011001", pass => true),
  (xin_0 => "001010101001111100", xin_1 => "000110010101000000", pass => true),
  (xin_0 => "001000100110000100", xin_1 => "000010010111110101", pass => false),
  (xin_0 => "001010011101010110", xin_1 => "001010000010101101", pass => false),
  (xin_0 => "001100100110101111", xin_1 => "000010011010101011", pass => true),
  (xin_0 => "000011110011100100", xin_1 => "001000101101111001", pass => false),
  (xin_0 => "001001110110010011", xin_1 => "000101101100011111", pass => true),
  (xin_0 => "001100101111110110", xin_1 => "001000001000101010", pass => false),
  (xin_0 => "000111011011000001", xin_1 => "000010011110100110", pass => false),
  (xin_0 => "001000001101110000", xin_1 => "000111011001110010", pass => true),
  (xin_0 => "001100001111001000", xin_1 => "000100100101010010", pass => true),
  (xin_0 => "000100100011101110", xin_1 => "000001111110011110", pass => true),
  (xin_0 => "001010110001100110", xin_1 => "000100010110100100", pass => true),
  (xin_0 => "001100011101100000", xin_1 => "000101110100111011", pass => false),
  (xin_0 => "000100011000101110", xin_1 => "001000000000111010", pass => false),
  (xin_0 => "000111011001000010", xin_1 => "001000001100101010", pass => true),
  (xin_0 => "000100001101100110", xin_1 => "000011000011001111", pass => true),
  (xin_0 => "001011110010000010", xin_1 => "001001111110111111", pass => false),
  (xin_0 => "000101011000111000", xin_1 => "000101001101010000", pass => true),
  (xin_0 => "001101000100010110", xin_1 => "000100000110111110", pass => true),
  (xin_0 => "001011011110011110", xin_1 => "001010001001010101", pass => false),
  (xin_0 => "000110111001001011", xin_1 => "000111101001000111", pass => true),
  (xin_0 => "001010001000000100", xin_1 => "001100000110001110", pass => false),
  (xin_0 => "001001000111110101", xin_1 => "000100010010100010", pass => true),
  (xin_0 => "000110011111111101", xin_1 => "000101100101001010", pass => true),
  (xin_0 => "001000010100101001", xin_1 => "000001010001011110", pass => false),
  (xin_0 => "001001110100011010", xin_1 => "001010110110000101", pass => false),
  (xin_0 => "001100011010000101", xin_1 => "001000000010001110", pass => false),
  (xin_0 => "000110101100011011", xin_1 => "000001100111101110", pass => false),
  (xin_0 => "001000100110011011", xin_1 => "000010110000010110", pass => false),
  (xin_0 => "000100111011011011", xin_1 => "000100110110110111", pass => true),
  (xin_0 => "000110010110001100", xin_1 => "001000110101100010", pass => false),
  (xin_0 => "001110101101000110", xin_1 => "000111011111101010", pass => false),
  (xin_0 => "000111011110010011", xin_1 => "000011111111110101", pass => false),
  (xin_0 => "001101000100111011", xin_1 => "001010110001000001", pass => true),
  (xin_0 => "001001001110111100", xin_1 => "000001111101010010", pass => false),
  (xin_0 => "000100101111110100", xin_1 => "000010010011100101", pass => true),
  (xin_0 => "001000000010011111", xin_1 => "000010000101011001", pass => false),
  (xin_0 => "000110101110011011", xin_1 => "000001110010001100", pass => false),
  (xin_0 => "000111001011010010", xin_1 => "001001100100001101", pass => false),
  (xin_0 => "000100100100001011", xin_1 => "000101011110010100", pass => true),
  (xin_0 => "000111111001001011", xin_1 => "000001100111010011", pass => false),
  (xin_0 => "000111011010110100", xin_1 => "000010100001101101", pass => false),
  (xin_0 => "000110101001101010", xin_1 => "001001110010100010", pass => false),
  (xin_0 => "000111110000001011", xin_1 => "000010010101100110", pass => false),
  (xin_0 => "000111010101011111", xin_1 => "000000111110000100", pass => false),
  (xin_0 => "000101001011111110", xin_1 => "000111101001110001", pass => false),
  (xin_0 => "000110101011001011", xin_1 => "000100010010000111", pass => true),
  (xin_0 => "001000010010110100", xin_1 => "000011000000011000", pass => false),
  (xin_0 => "001101011111010010", xin_1 => "000011011101101110", pass => true),
  (xin_0 => "001010011100010011", xin_1 => "001000011001101000", pass => false),
  (xin_0 => "001000111001001010", xin_1 => "000010110000110110", pass => false),
  (xin_0 => "000110110010001101", xin_1 => "000110000111111100", pass => true),
  (xin_0 => "001111001110111000", xin_1 => "001001000010101010", pass => true),
  (xin_0 => "000111010000101001", xin_1 => "000110100000110011", pass => true),
  (xin_0 => "001100010111100011", xin_1 => "000110001000000011", pass => false),
  (xin_0 => "001000110010101111", xin_1 => "000010010100100111", pass => false),
  (xin_0 => "000100110000000001", xin_1 => "000111010111111111", pass => false),
  (xin_0 => "001011010100101100", xin_1 => "001000110010111100", pass => false),
  (xin_0 => "000101111111000011", xin_1 => "000100110011010010", pass => true),
  (xin_0 => "000100100011000110", xin_1 => "001000001110110111", pass => false),
  (xin_0 => "001100010100001111", xin_1 => "000010111100011000", pass => true),
  (xin_0 => "001111111111110100", xin_1 => "001010001101001110", pass => true),
  (xin_0 => "000111001111011010", xin_1 => "000010111100110100", pass => false),
  (xin_0 => "001011111100100110", xin_1 => "000111000100111101", pass => false),
  (xin_0 => "001001000101000001", xin_1 => "000001111111110011", pass => false),
  (xin_0 => "001001011000011100", xin_1 => "001010000100010101", pass => false),
  (xin_0 => "001100101100100010", xin_1 => "001000001011110011", pass => false),
  (xin_0 => "000101111011101110", xin_1 => "000010111101110000", pass => false),
  (xin_0 => "001001001101100100", xin_1 => "000010111000101010", pass => false),
  (xin_0 => "000011111011000101", xin_1 => "000111000000000001", pass => false),
  (xin_0 => "001011001010010011", xin_1 => "000110100110110111", pass => true),
  (xin_0 => "001000100001100101", xin_1 => "001011000110011000", pass => false),
  (xin_0 => "001011101011001011", xin_1 => "000101001010001110", pass => true),
  (xin_0 => "001001001101011011", xin_1 => "000010100000111111", pass => false),
  (xin_0 => "001001101111010000", xin_1 => "000010010100101001", pass => false),
  (xin_0 => "001001100011111101", xin_1 => "001100110111011000", pass => false),
  (xin_0 => "000011110000010011", xin_1 => "000011010100111111", pass => true),
  (xin_0 => "000110000010100111", xin_1 => "000010010100011110", pass => false),
  (xin_0 => "000110011110011101", xin_1 => "001010100111000111", pass => false),
  (xin_0 => "001011011010000000", xin_1 => "001010011110000110", pass => false),
  (xin_0 => "000111001111001000", xin_1 => "000001011011111000", pass => false),
  (xin_0 => "001000110100000100", xin_1 => "001010110110001000", pass => false),
  (xin_0 => "001001110100011101", xin_1 => "001010110001001110", pass => false),
  (xin_0 => "001000001101000010", xin_1 => "001010010010110000", pass => false),
  (xin_0 => "001101010111100010", xin_1 => "000011101001001111", pass => true),
  (xin_0 => "001001111000011100", xin_1 => "000111011011000111", pass => true),
  (xin_0 => "000100010101001000", xin_1 => "000001110111010101", pass => true),
  (xin_0 => "000111000001101100", xin_1 => "000011000100011110", pass => false),
  (xin_0 => "000111111110110001", xin_1 => "000110110010000010", pass => true),
  (xin_0 => "001000100000001011", xin_1 => "000011000101110111", pass => false),
  (xin_0 => "001010001111010011", xin_1 => "001100010010010010", pass => false),
  (xin_0 => "000101001011000101", xin_1 => "000010101011101110", pass => true),
  (xin_0 => "001011011001010010", xin_1 => "001000001001111101", pass => false),
  (xin_0 => "001010001111010110", xin_1 => "001001101101000011", pass => false),
  (xin_0 => "000111101111011110", xin_1 => "000010011010000101", pass => false),
  (xin_0 => "000101011010010101", xin_1 => "000100001010010100", pass => true),
  (xin_0 => "001000111000111001", xin_1 => "000101100111001011", pass => true),
  (xin_0 => "000101111110111111", xin_1 => "001010110111100110", pass => false),
  (xin_0 => "001000110101011110", xin_1 => "001100100101011111", pass => false),
  (xin_0 => "001010101101000000", xin_1 => "001001010110011100", pass => false),
  (xin_0 => "001001101010010011", xin_1 => "001010100011000100", pass => false),
  (xin_0 => "001100010111101100", xin_1 => "001000100011100111", pass => false),
  (xin_0 => "001100110111010010", xin_1 => "000101101100001100", pass => false),
  (xin_0 => "001001010011110110", xin_1 => "000001010011011010", pass => false),
  (xin_0 => "000110000011001010", xin_1 => "000011100010011011", pass => false),
  (xin_0 => "000110011111011101", xin_1 => "001001001001110111", pass => false),
  (xin_0 => "001110111101100000", xin_1 => "001001111010011101", pass => true),
  (xin_0 => "001000000000101001", xin_1 => "000111011010000100", pass => true),
  (xin_0 => "000101011010001001", xin_1 => "000101110111100000", pass => true),
  (xin_0 => "001011001101011111", xin_1 => "000011110000000110", pass => true),
  (xin_0 => "001001001110111101", xin_1 => "000101100010101101", pass => true),
  (xin_0 => "001010111000101001", xin_1 => "000011001001110111", pass => true),
  (xin_0 => "001010100000010111", xin_1 => "001001000001110001", pass => false),
  (xin_0 => "001100100100101001", xin_1 => "001000101001000001", pass => false),
  (xin_0 => "000110111100000011", xin_1 => "001001100001100000", pass => false),
  (xin_0 => "001101010110111010", xin_1 => "000111011110001101", pass => false),
  (xin_0 => "001001010101101101", xin_1 => "000100100000000101", pass => true),
  (xin_0 => "001000111110000011", xin_1 => "000010110000000000", pass => false),
  (xin_0 => "001000100101010001", xin_1 => "000010110000100101", pass => false),
  (xin_0 => "000011100101101010", xin_1 => "000111111000100011", pass => false),
  (xin_0 => "000101100111000010", xin_1 => "001000000000110101", pass => false),
  (xin_0 => "000110000000011011", xin_1 => "000101110010001001", pass => true),
  (xin_0 => "001101100010110110", xin_1 => "000100110011100011", pass => false),
  (xin_0 => "000111101000010101", xin_1 => "000101001111111111", pass => true),
  (xin_0 => "001101011100001011", xin_1 => "000111101100010001", pass => false),
  (xin_0 => "001000111011101101", xin_1 => "000010101110100111", pass => false),
  (xin_0 => "001100100000100001", xin_1 => "111111100010101110", pass => true),
  (xin_0 => "001100011010011010", xin_1 => "000101010000100001", pass => true),
  (xin_0 => "000011101011111111", xin_1 => "000100000101011010", pass => true),
  (xin_0 => "000111110000101010", xin_1 => "000100001000100010", pass => false),
  (xin_0 => "000110010001010000", xin_1 => "001001000000101101", pass => false),
  (xin_0 => "001100000011000000", xin_1 => "001000010000011100", pass => false),
  (xin_0 => "000111000111000110", xin_1 => "001011011101011000", pass => false),
  (xin_0 => "000110100100010001", xin_1 => "000100110010111000", pass => true),
  (xin_0 => "000011111000001100", xin_1 => "001000011010111110", pass => false),
  (xin_0 => "000101101111000101", xin_1 => "001001100101001011", pass => false),
  (xin_0 => "001011010110111110", xin_1 => "001000010101010000", pass => false),
  (xin_0 => "001000010110001010", xin_1 => "000111010001100111", pass => true),
  (xin_0 => "000110100011011110", xin_1 => "000011101011010001", pass => false),
  (xin_0 => "001010000100111110", xin_1 => "000111101100110001", pass => true),
  (xin_0 => "001100000010111011", xin_1 => "000111111101111101", pass => false),
  (xin_0 => "000101001010010101", xin_1 => "000110011100010101", pass => true),
  (xin_0 => "000101011001010110", xin_1 => "000011110001110010", pass => true),
  (xin_0 => "000110000001000001", xin_1 => "000101000111111010", pass => true),
  (xin_0 => "001010010101111011", xin_1 => "001010101101110101", pass => false),
  (xin_0 => "001100101000011111", xin_1 => "000111100010101111", pass => false),
  (xin_0 => "001001000000100110", xin_1 => "000010110011100011", pass => false),
  (xin_0 => "000011010101001011", xin_1 => "000001010101011011", pass => true),
  (xin_0 => "000110100110100100", xin_1 => "000010000111111000", pass => false),
  (xin_0 => "001001110111000111", xin_1 => "000110110011010001", pass => true),
  (xin_0 => "001010000001111000", xin_1 => "000010011111110101", pass => false),
  (xin_0 => "001011000000001010", xin_1 => "001001000110111011", pass => false),
  (xin_0 => "001001010111001010", xin_1 => "000110100000111111", pass => true),
  (xin_0 => "000100110011010010", xin_1 => "000010101000100011", pass => true),
  (xin_0 => "001001101111011011", xin_1 => "000010110100000101", pass => false),
  (xin_0 => "001000111101000110", xin_1 => "000111000101011101", pass => true),
  (xin_0 => "001010101001101010", xin_1 => "000101011001011101", pass => true),
  (xin_0 => "001011010110011011", xin_1 => "001000100001011100", pass => false),
  (xin_0 => "001000010100011011", xin_1 => "000110100111011111", pass => true),
  (xin_0 => "001011011000000101", xin_1 => "001000110011110011", pass => false),
  (xin_0 => "001001110001000101", xin_1 => "000101000000110010", pass => true),
  (xin_0 => "000101011111110111", xin_1 => "000100100111100011", pass => true),
  (xin_0 => "001001110110110101", xin_1 => "000010011111111010", pass => false),
  (xin_0 => "000110100110010010", xin_1 => "000010011110100011", pass => false),
  (xin_0 => "000111111101110010", xin_1 => "000110000111100110", pass => true),
  (xin_0 => "000100011111100001", xin_1 => "001000001011100111", pass => false),
  (xin_0 => "000110000010011110", xin_1 => "000101111100111001", pass => true),
  (xin_0 => "001001111000100100", xin_1 => "000111001000110000", pass => true),
  (xin_0 => "000111100010100010", xin_1 => "000010010000011100", pass => false),
  (xin_0 => "001000000010000110", xin_1 => "000111001100010001", pass => true),
  (xin_0 => "001000101100110011", xin_1 => "000010111101101110", pass => false),
  (xin_0 => "001101000001011000", xin_1 => "000111010111111101", pass => false),
  (xin_0 => "001010011001111100", xin_1 => "000110011001010100", pass => true),
  (xin_0 => "001001000001010111", xin_1 => "000101101011100100", pass => true),
  (xin_0 => "000100101010000011", xin_1 => "000100001001111000", pass => true),
  (xin_0 => "001011001111111001", xin_1 => "001001001110101110", pass => false),
  (xin_0 => "001011011100010101", xin_1 => "000011010101011010", pass => true),
  (xin_0 => "000111010110110101", xin_1 => "000111000110100000", pass => true),
  (xin_0 => "001110100101010101", xin_1 => "000100010000001010", pass => false),
  (xin_0 => "001101100100001111", xin_1 => "000101111001000010", pass => false),
  (xin_0 => "001011000100101000", xin_1 => "001010001100111001", pass => false),
  (xin_0 => "001001111111010010", xin_1 => "001000001100011000", pass => false),
  (xin_0 => "000011110110101010", xin_1 => "000010001011011001", pass => true),
  (xin_0 => "001001000111010111", xin_1 => "001011111011010111", pass => false),
  (xin_0 => "000110001001010011", xin_1 => "001001010101110110", pass => false),
  (xin_0 => "000101001001111100", xin_1 => "000010110111000010", pass => true),
  (xin_0 => "001100010001101011", xin_1 => "000111111100011001", pass => false),
  (xin_0 => "000111001001000100", xin_1 => "000010110000011100", pass => false),
  (xin_0 => "001100110001011111", xin_1 => "000110111000111010", pass => false),
  (xin_0 => "010000000001100110", xin_1 => "001010011001010000", pass => true),
  (xin_0 => "001110100101011001", xin_1 => "001010000001101011", pass => true),
  (xin_0 => "000111100101101111", xin_1 => "000011011011110100", pass => false),
  (xin_0 => "001100001011110100", xin_1 => "000100110111100100", pass => true),
  (xin_0 => "000011110100110101", xin_1 => "000100011011010111", pass => true),
  (xin_0 => "001010000101111011", xin_1 => "001011001101001100", pass => false),
  (xin_0 => "001010011011101100", xin_1 => "000011111000001100", pass => true),
  (xin_0 => "001101110001100000", xin_1 => "000101000011110110", pass => false),
  (xin_0 => "001000010000000110", xin_1 => "000001110000101000", pass => false),
  (xin_0 => "000110111001001101", xin_1 => "001001001001010101", pass => false),
  (xin_0 => "001011101100110111", xin_1 => "001010100001000101", pass => false),
  (xin_0 => "001001001110000011", xin_1 => "000101110000100110", pass => true),
  (xin_0 => "000111011100101000", xin_1 => "001010010110001011", pass => false),
  (xin_0 => "000100000110111011", xin_1 => "000101011010110001", pass => true),
  (xin_0 => "000111001001001001", xin_1 => "001001101011100111", pass => false),
  (xin_0 => "001100010000100110", xin_1 => "000101010110111011", pass => true),
  (xin_0 => "001110100000001101", xin_1 => "000110010110111001", pass => false),
  (xin_0 => "000110111101100100", xin_1 => "000100110101100001", pass => true),
  (xin_0 => "001001001111111110", xin_1 => "000011000101110001", pass => false),
  (xin_0 => "001011001110101100", xin_1 => "001001000110011101", pass => false),
  (xin_0 => "001001001000010001", xin_1 => "000010011111000100", pass => false),
  (xin_0 => "000111001001000000", xin_1 => "000010101000110011", pass => false),
  (xin_0 => "001010011010000100", xin_1 => "000100100110001101", pass => true),
  (xin_0 => "001001000110111111", xin_1 => "000011001001011010", pass => false),
  (xin_0 => "001011110010101010", xin_1 => "000110000110000001", pass => true),
  (xin_0 => "001000111000100110", xin_1 => "000110001110101001", pass => true),
  (xin_0 => "001010001110101001", xin_1 => "000111011100000110", pass => true),
  (xin_0 => "000110111001010000", xin_1 => "000111101001000111", pass => true),
  (xin_0 => "001100100100001011", xin_1 => "000101110111100010", pass => false),
  (xin_0 => "001010010101011101", xin_1 => "001011110001111011", pass => false),
  (xin_0 => "001011110110000000", xin_1 => "000111010110100101", pass => false),
  (xin_0 => "001101000100110100", xin_1 => "000010111000100111", pass => true),
  (xin_0 => "001011111001111111", xin_1 => "000100100011101110", pass => true),
  (xin_0 => "000110001101100100", xin_1 => "001001010100010100", pass => false),
  (xin_0 => "000011110101011100", xin_1 => "000011011011000001", pass => true),
  (xin_0 => "001100110001000100", xin_1 => "000100010110110001", pass => true),
  (xin_0 => "000110101111110100", xin_1 => "000111010111001011", pass => true),
  (xin_0 => "001100100011101011", xin_1 => "001000000100110111", pass => false),
  (xin_0 => "001100111100000100", xin_1 => "000010000101101101", pass => true),
  (xin_0 => "000100010100010000", xin_1 => "001000001001011111", pass => false),
  (xin_0 => "000111000111100001", xin_1 => "001011001110110010", pass => false),
  (xin_0 => "000100110000111001", xin_1 => "000101100110111111", pass => true),
  (xin_0 => "001000000101101100", xin_1 => "000010011010010101", pass => false),
  (xin_0 => "001000010000101111", xin_1 => "000010101011010111", pass => false),
  (xin_0 => "001011011111110001", xin_1 => "000011101000000001", pass => true),
  (xin_0 => "000110101011110010", xin_1 => "000010001011010010", pass => false),
  (xin_0 => "000110101001100011", xin_1 => "000001111001010100", pass => false),
  (xin_0 => "000100110111101101", xin_1 => "000011001000000100", pass => true),
  (xin_0 => "000110000101111111", xin_1 => "000011111111101001", pass => true),
  (xin_0 => "001101010101111100", xin_1 => "000101001001011111", pass => false),
  (xin_0 => "001000111010010100", xin_1 => "000010101110011111", pass => false),
  (xin_0 => "000100110110000100", xin_1 => "000010010100101011", pass => true),
  (xin_0 => "001101001011010110", xin_1 => "000110010101110100", pass => false),
  (xin_0 => "001010111001011101", xin_1 => "000110110001101110", pass => true),
  (xin_0 => "001000100011111110", xin_1 => "000110101001000011", pass => true),
  (xin_0 => "001000000001101111", xin_1 => "001000011000001001", pass => true),
  (xin_0 => "001001011110010000", xin_1 => "001011111001101111", pass => false),
  (xin_0 => "001100000011101100", xin_1 => "000111100111011011", pass => false),
  (xin_0 => "000100100100011111", xin_1 => "000101011010000000", pass => true),
  (xin_0 => "001000011110010100", xin_1 => "000011001110110001", pass => false),
  (xin_0 => "001000010101011000", xin_1 => "001011100100001010", pass => false),
  (xin_0 => "001010101010010110", xin_1 => "000011110011110001", pass => true),
  (xin_0 => "000111110110101101", xin_1 => "000001010111011010", pass => false),
  (xin_0 => "001011101101100001", xin_1 => "001000000110010100", pass => false),
  (xin_0 => "001000011010010101", xin_1 => "000010000001100110", pass => false),
  (xin_0 => "000100010111101011", xin_1 => "000010011010011111", pass => true),
  (xin_0 => "000110110010000100", xin_1 => "000110010000100001", pass => true),
  (xin_0 => "000100000001010000", xin_1 => "000010101101001111", pass => true),
  (xin_0 => "001010011100001110", xin_1 => "001010110001011111", pass => false),
  (xin_0 => "001001100110111101", xin_1 => "000010000001001101", pass => false),
  (xin_0 => "001010101111011101", xin_1 => "001001100101110000", pass => false),
  (xin_0 => "001010010100100100", xin_1 => "000111000110111000", pass => true),
  (xin_0 => "000101011000001110", xin_1 => "000010101110110110", pass => true),
  (xin_0 => "001100001011111010", xin_1 => "001001010010100010", pass => false),
  (xin_0 => "001010111011000101", xin_1 => "001000011110010111", pass => false),
  (xin_0 => "001011000110000110", xin_1 => "001000010001100100", pass => false),
  (xin_0 => "000111110011100000", xin_1 => "000001110100001110", pass => false),
  (xin_0 => "001000110100001011", xin_1 => "000010011110000100", pass => false),
  (xin_0 => "000100110001000011", xin_1 => "000110000000000011", pass => true),
  (xin_0 => "001111101011110011", xin_1 => "001010010000000110", pass => true),
  (xin_0 => "001100000000011100", xin_1 => "000101001000001001", pass => true),
  (xin_0 => "001011111111101000", xin_1 => "000011000001110100", pass => true),
  (xin_0 => "001001001010101011", xin_1 => "000110100110101001", pass => true),
  (xin_0 => "001110000101101101", xin_1 => "000110100011101110", pass => false),
  (xin_0 => "001001101010110100", xin_1 => "000111011110010100", pass => true),
  (xin_0 => "001001010110111111", xin_1 => "001010000000111111", pass => false),
  (xin_0 => "000100011010011000", xin_1 => "000101100110101110", pass => true),
  (xin_0 => "001110011011100100", xin_1 => "001010010011111001", pass => true),
  (xin_0 => "000111100000011100", xin_1 => "000101011111101101", pass => true),
  (xin_0 => "001010010011001100", xin_1 => "000010011001110101", pass => false),
  (xin_0 => "000110000100101110", xin_1 => "001001101100101010", pass => false),
  (xin_0 => "000110110001001010", xin_1 => "001001110110010011", pass => false),
  (xin_0 => "001001010110110100", xin_1 => "000011111010011010", pass => false),
  (xin_0 => "000111001011010111", xin_1 => "001000100101011000", pass => true),
  (xin_0 => "001001011010011010", xin_1 => "001000000000100001", pass => true),
  (xin_0 => "000100111101110011", xin_1 => "001000010010100000", pass => false),
  (xin_0 => "001010011110011110", xin_1 => "001010101101100100", pass => false),
  (xin_0 => "000111001011111101", xin_1 => "000101010011000011", pass => true),
  (xin_0 => "001100001111111000", xin_1 => "001000001100010110", pass => false),
  (xin_0 => "000101011101110110", xin_1 => "001001000011111000", pass => false),
  (xin_0 => "000110010001000100", xin_1 => "000100111111101001", pass => true),
  (xin_0 => "001010110111100111", xin_1 => "000101100111110110", pass => true),
  (xin_0 => "000101001110111011", xin_1 => "000101011100010000", pass => true),
  (xin_0 => "001001001101111000", xin_1 => "000001111111001100", pass => false),
  (xin_0 => "001001110001011010", xin_1 => "000111011011010001", pass => true),
  (xin_0 => "000100001100111110", xin_1 => "000101110111000100", pass => true),
  (xin_0 => "001011110001101100", xin_1 => "000111110010001100", pass => false),
  (xin_0 => "001010111101110111", xin_1 => "001000001101010010", pass => false),
  (xin_0 => "000111100000110010", xin_1 => "000010010011000001", pass => false),
  (xin_0 => "001001000001011000", xin_1 => "000010111110111101", pass => false),
  (xin_0 => "001001010101011100", xin_1 => "001100010011001000", pass => false),
  (xin_0 => "001001110100110011", xin_1 => "000010101010100000", pass => false),
  (xin_0 => "001000101111100101", xin_1 => "000100111011010001", pass => true),
  (xin_0 => "000100100001010010", xin_1 => "001000001110100101", pass => false),
  (xin_0 => "001101010000110000", xin_1 => "000101110000010001", pass => false),
  (xin_0 => "001110110000011011", xin_1 => "001010001000010101", pass => true),
  (xin_0 => "000111110110000100", xin_1 => "000010011001110011", pass => false),
  (xin_0 => "000111101001001101", xin_1 => "000111110100100011", pass => true),
  (xin_0 => "000110111000111000", xin_1 => "000010111000111011", pass => false),
  (xin_0 => "001000100001101100", xin_1 => "001011110110111100", pass => false),
  (xin_0 => "000110100000110001", xin_1 => "000010111100100000", pass => false),
  (xin_0 => "000110100101111011", xin_1 => "000111001111100000", pass => true),
  (xin_0 => "000110010011011111", xin_1 => "001001011110000101", pass => false),
  (xin_0 => "001001010110010101", xin_1 => "000011100110110101", pass => false),
  (xin_0 => "001000011001010011", xin_1 => "000101010110011101", pass => true),
  (xin_0 => "000011010101010110", xin_1 => "001000000010111011", pass => false),
  (xin_0 => "000100111110100011", xin_1 => "000011011110101110", pass => true),
  (xin_0 => "001100000111111010", xin_1 => "000100010001011100", pass => true),
  (xin_0 => "001001110001100101", xin_1 => "001011111000100011", pass => false),
  (xin_0 => "001000101010010101", xin_1 => "000011111001101101", pass => false),
  (xin_0 => "001011100110010111", xin_1 => "000101010000101111", pass => true),
  (xin_0 => "001000001011010101", xin_1 => "001000100000100010", pass => true),
  (xin_0 => "001100100110000000", xin_1 => "111110111110011001", pass => true),
  (xin_0 => "001100010111011111", xin_1 => "000101001101011100", pass => true),
  (xin_0 => "001011010111101111", xin_1 => "001001111110111110", pass => false),
  (xin_0 => "000111000111011111", xin_1 => "000011010010001000", pass => false),
  (xin_0 => "000011110000011000", xin_1 => "000110000000011010", pass => true),
  (xin_0 => "001110110111001110", xin_1 => "000100110100101111", pass => false),
  (xin_0 => "001100011000101110", xin_1 => "001010110000000001", pass => false),
  (xin_0 => "001000110111010110", xin_1 => "000010111001101111", pass => false),
  (xin_0 => "001011011011101110", xin_1 => "001000010000101011", pass => false),
  (xin_0 => "001001101111010001", xin_1 => "000110011010001001", pass => true),
  (xin_0 => "001001111011000001", xin_1 => "001001011001101010", pass => false),
  (xin_0 => "000110101111100010", xin_1 => "000100011111000101", pass => true),
  (xin_0 => "001000111000010001", xin_1 => "000010010001101110", pass => false),
  (xin_0 => "001101000111111001", xin_1 => "000111000100010000", pass => false),
  (xin_0 => "001001101100111001", xin_1 => "000111101100010011", pass => true),
  (xin_0 => "000110011011111001", xin_1 => "001010011011000100", pass => false),
  (xin_0 => "000101110000011011", xin_1 => "000111001101001001", pass => true),
  (xin_0 => "000101000100011000", xin_1 => "000011000010110001", pass => true),
  (xin_0 => "000110000111010100", xin_1 => "000001101101011000", pass => false),
  (xin_0 => "001001101101010010", xin_1 => "000100100101011111", pass => true),
  (xin_0 => "000011110011011011", xin_1 => "000101000100111110", pass => true),
  (xin_0 => "001110111011100010", xin_1 => "000100110000111000", pass => false),
  (xin_0 => "001001100001110011", xin_1 => "000010100111011001", pass => false),
  (xin_0 => "000101110110010100", xin_1 => "000100010110101101", pass => true),
  (xin_0 => "001101010000111011", xin_1 => "000110001101000011", pass => false),
  (xin_0 => "000111111000101000", xin_1 => "001000010101000111", pass => true),
  (xin_0 => "001100011101010010", xin_1 => "001010000111110011", pass => false),
  (xin_0 => "001001111101010101", xin_1 => "000101011111100000", pass => true),
  (xin_0 => "001010001110101001", xin_1 => "001001101111101001", pass => false),
  (xin_0 => "000111000001110000", xin_1 => "001001111101011000", pass => false),
  (xin_0 => "000111011110001101", xin_1 => "001010110001101011", pass => false),
  (xin_0 => "000110011000110001", xin_1 => "000010010111110110", pass => false),
  (xin_0 => "001100111100001111", xin_1 => "001010000010000000", pass => true),
  (xin_0 => "001000011001010110", xin_1 => "001011010000110111", pass => false),
  (xin_0 => "000101111110100001", xin_1 => "001010001101000100", pass => false),
  (xin_0 => "000111100101010100", xin_1 => "000110011111000110", pass => true),
  (xin_0 => "000101101010110100", xin_1 => "001001000011000100", pass => false),
  (xin_0 => "001010001000000101", xin_1 => "000100100010100101", pass => true),
  (xin_0 => "001110110110000101", xin_1 => "000100111011100001", pass => false),
  (xin_0 => "000110101111101100", xin_1 => "000010110111001001", pass => false),
  (xin_0 => "000111011110111110", xin_1 => "001000010100101111", pass => true),
  (xin_0 => "000101010100011000", xin_1 => "000111101011101101", pass => false),
  (xin_0 => "000110100101000100", xin_1 => "000010100011101010", pass => false),
  (xin_0 => "000110010011000110", xin_1 => "000111011011110100", pass => true),
  (xin_0 => "000101100000100001", xin_1 => "001001101011101111", pass => false),
  (xin_0 => "000111011101010101", xin_1 => "000011011000101101", pass => false),
  (xin_0 => "001010110000111011", xin_1 => "001011010011011111", pass => false),
  (xin_0 => "001100011011011001", xin_1 => "000011111011111110", pass => true),
  (xin_0 => "001100111110110110", xin_1 => "000101100100000101", pass => false),
  (xin_0 => "001000100101001010", xin_1 => "000110000010101101", pass => true),
  (xin_0 => "000111000100000010", xin_1 => "000010110111101110", pass => false),
  (xin_0 => "001001010000001101", xin_1 => "000011000011011010", pass => false),
  (xin_0 => "000111001010101000", xin_1 => "001011001000101111", pass => false),
  (xin_0 => "001100100111001011", xin_1 => "000101011101110110", pass => false),
  (xin_0 => "000100110100110011", xin_1 => "001000110000000000", pass => false),
  (xin_0 => "000100101101000101", xin_1 => "000011101111101010", pass => true),
  (xin_0 => "001100110001100000", xin_1 => "000110100000100111", pass => false),
  (xin_0 => "000111011001101001", xin_1 => "000011110000001101", pass => false),
  (xin_0 => "000111110100100000", xin_1 => "001001010110101110", pass => false),
  (xin_0 => "000110010101101011", xin_1 => "000101001000100010", pass => true),
  (xin_0 => "001000111111010100", xin_1 => "000100001101010001", pass => false),
  (xin_0 => "001101001110011001", xin_1 => "000001110101101011", pass => true),
  (xin_0 => "000111100100011101", xin_1 => "001000010010000101", pass => true),
  (xin_0 => "000111100100001100", xin_1 => "000110011100100011", pass => true),
  (xin_0 => "001010011100010100", xin_1 => "001010000101011110", pass => false),
  (xin_0 => "001100000000100010", xin_1 => "000111011110001110", pass => false),
  (xin_0 => "001010011110101111", xin_1 => "000010110011001100", pass => false),
  (xin_0 => "000111111000100101", xin_1 => "000010110000011110", pass => false),
  (xin_0 => "001100101011111110", xin_1 => "000111000101100110", pass => false),
  (xin_0 => "000101111100110010", xin_1 => "000101110101001001", pass => true),
  (xin_0 => "000101101100100001", xin_1 => "001001100101000100", pass => false),
  (xin_0 => "001000011010110011", xin_1 => "000001111101101000", pass => false),
  (xin_0 => "001011101001100111", xin_1 => "001000100110111111", pass => false),
  (xin_0 => "001001011100010000", xin_1 => "001011011010000011", pass => false),
  (xin_0 => "001000111000110010", xin_1 => "000110101110010100", pass => true),
  (xin_0 => "000101001010110001", xin_1 => "000110100101011011", pass => true),
  (xin_0 => "001100110110010111", xin_1 => "001010100110100011", pass => true),
  (xin_0 => "001110000000100110", xin_1 => "000101110010110100", pass => false),
  (xin_0 => "000101010111000010", xin_1 => "000100000010100011", pass => true),
  (xin_0 => "001000111000011011", xin_1 => "000001101011100111", pass => false),
  (xin_0 => "001010011000110011", xin_1 => "001010111010110101", pass => false),
  (xin_0 => "001010100011000111", xin_1 => "001010101101110111", pass => false),
  (xin_0 => "001010001100000001", xin_1 => "000110110100010001", pass => true),
  (xin_0 => "001101101110000001", xin_1 => "000100011000110010", pass => false),
  (xin_0 => "001010100011101001", xin_1 => "000011101111101001", pass => true),
  (xin_0 => "000101111100110010", xin_1 => "001010010001110000", pass => false),
  (xin_0 => "001001110011110010", xin_1 => "000010000101001110", pass => false),
  (xin_0 => "001101000110100110", xin_1 => "000101000111010011", pass => false),
  (xin_0 => "001010001111101010", xin_1 => "000010111110000101", pass => false),
  (xin_0 => "000110110100111100", xin_1 => "001000111010000011", pass => false),
  (xin_0 => "001010001000101111", xin_1 => "000110010010000011", pass => true),
  (xin_0 => "001001001001111111", xin_1 => "001011011001111000", pass => false),
  (xin_0 => "001100011011100101", xin_1 => "000011010110111010", pass => true),
  (xin_0 => "001001110100111001", xin_1 => "000011011010000001", pass => false),
  (xin_0 => "000111100010101000", xin_1 => "000010110010010000", pass => false),
  (xin_0 => "000110011110001011", xin_1 => "000010010000010111", pass => false),
  (xin_0 => "001011010001111110", xin_1 => "001010010110000101", pass => false),
  (xin_0 => "001000011101010010", xin_1 => "000110010000100110", pass => true),
  (xin_0 => "000111110111010101", xin_1 => "000011010000111010", pass => false),
  (xin_0 => "000110100001111100", xin_1 => "000100010000001000", pass => true),
  (xin_0 => "001011000101101100", xin_1 => "000101101010111100", pass => true),
  (xin_0 => "000101011101001101", xin_1 => "001010000101001111", pass => false),
  (xin_0 => "000101101101000111", xin_1 => "000010100101100101", pass => false),
  (xin_0 => "001010000100000000", xin_1 => "000011001110100000", pass => false),
  (xin_0 => "001011000111001010", xin_1 => "000111010101101111", pass => false),
  (xin_0 => "000100000000111000", xin_1 => "000111100000101111", pass => false),
  (xin_0 => "000100011110000100", xin_1 => "000100010111110110", pass => true),
  (xin_0 => "001000111101110110", xin_1 => "001010101100000011", pass => false),
  (xin_0 => "001100111011000111", xin_1 => "000011110010110101", pass => true),
  (xin_0 => "000110011010011000", xin_1 => "000111000001110011", pass => true),
  (xin_0 => "000101011111011000", xin_1 => "001000001110110000", pass => false),
  (xin_0 => "001010100011011000", xin_1 => "000101011111000111", pass => true),
  (xin_0 => "001010111001110110", xin_1 => "000110110000000000", pass => true),
  (xin_0 => "001010001000011000", xin_1 => "000100000101000000", pass => true),
  (xin_0 => "000110001010110010", xin_1 => "001000100001011010", pass => false),
  (xin_0 => "000101101101111011", xin_1 => "000111111110101110", pass => false),
  (xin_0 => "000011101011110010", xin_1 => "000011101001101101", pass => true),
  (xin_0 => "001010011100011000", xin_1 => "001010110111000111", pass => false),
  (xin_0 => "000111100001110110", xin_1 => "000110100110101101", pass => true),
  (xin_0 => "001010111100111011", xin_1 => "001011000000000000", pass => false),
  (xin_0 => "000100111101011110", xin_1 => "000101010000010001", pass => true),
  (xin_0 => "001110101010011110", xin_1 => "000011111000010111", pass => false),
  (xin_0 => "001001011011010010", xin_1 => "000010001110101111", pass => false),
  (xin_0 => "001101010110100000", xin_1 => "000010001010000100", pass => true),
  (xin_0 => "000111110000110010", xin_1 => "000010010001111010", pass => false),
  (xin_0 => "001001011101000010", xin_1 => "000100111011010001", pass => true),
  (xin_0 => "001000010001001111", xin_1 => "001010100110011100", pass => false),
  (xin_0 => "001011111111011011", xin_1 => "000111011011101111", pass => false),
  (xin_0 => "010000000110001110", xin_1 => "001001100111111111", pass => true),
  (xin_0 => "001011010110001101", xin_1 => "001010100010100101", pass => false),
  (xin_0 => "000111011000111110", xin_1 => "000010000000000011", pass => false),
  (xin_0 => "000100100001011001", xin_1 => "000111011010011100", pass => false),
  (xin_0 => "000101111101010111", xin_1 => "000010111010000100", pass => false),
  (xin_0 => "001010100011011001", xin_1 => "001001000101110001", pass => false),
  (xin_0 => "000110001111100001", xin_1 => "001011101110110001", pass => false),
  (xin_0 => "000011010101010111", xin_1 => "000101011001100000", pass => true),
  (xin_0 => "001100100010110110", xin_1 => "001000101011111101", pass => false),
  (xin_0 => "000111011010010001", xin_1 => "000010101011001001", pass => false),
  (xin_0 => "001001011010001010", xin_1 => "000100001111101110", pass => true),
  (xin_0 => "000100101011011100", xin_1 => "001000011110011110", pass => false),
  (xin_0 => "000101111100110101", xin_1 => "001000000111011011", pass => false),
  (xin_0 => "001100110101111001", xin_1 => "000000101111100000", pass => true),
  (xin_0 => "000011010001101110", xin_1 => "000100111000101010", pass => true),
  (xin_0 => "001001010010011001", xin_1 => "000100111000010100", pass => true),
  (xin_0 => "000100000100000010", xin_1 => "000100100101001011", pass => true),
  (xin_0 => "000101110001010111", xin_1 => "000010011101000101", pass => false),
  (xin_0 => "001000010101100111", xin_1 => "000010101000111110", pass => false),
  (xin_0 => "000011110010011001", xin_1 => "000100101111000010", pass => true),
  (xin_0 => "001000000100110110", xin_1 => "000011100010101110", pass => false),
  (xin_0 => "000101110001100100", xin_1 => "001000011101111110", pass => false),
  (xin_0 => "000101111110111111", xin_1 => "001000110011101110", pass => false),
  (xin_0 => "001010100100011000", xin_1 => "001010011011000011", pass => false),
  (xin_0 => "000101110101100000", xin_1 => "001010001100101101", pass => false),
  (xin_0 => "001001000011010111", xin_1 => "000010101001001000", pass => false),
  (xin_0 => "000111110111000011", xin_1 => "001000000100101101", pass => true),
  (xin_0 => "001110001100101010", xin_1 => "000101100100001111", pass => false),
  (xin_0 => "001001100010011010", xin_1 => "000010101010010110", pass => false),
  (xin_0 => "000100000101011110", xin_1 => "000111011011111010", pass => false),
  (xin_0 => "001001110011101110", xin_1 => "000101011001010111", pass => true),
  (xin_0 => "001000010000010010", xin_1 => "001000100101001100", pass => true),
  (xin_0 => "001010111111101001", xin_1 => "000011011101100111", pass => true),
  (xin_0 => "001000001001111010", xin_1 => "000010100110101001", pass => false),
  (xin_0 => "000011110011000100", xin_1 => "000001101100110010", pass => true),
  (xin_0 => "000111001000100001", xin_1 => "000101011010100110", pass => true),
  (xin_0 => "000111001111100110", xin_1 => "000010011110100100", pass => false),
  (xin_0 => "001010010110110100", xin_1 => "000010010001101011", pass => false),
  (xin_0 => "000101000000100010", xin_1 => "000101001111100010", pass => true),
  (xin_0 => "000111100110011000", xin_1 => "000011010110110010", pass => false),
  (xin_0 => "001001111000110110", xin_1 => "000011110011101000", pass => true),
  (xin_0 => "001101101001001101", xin_1 => "000101110101001011", pass => false),
  (xin_0 => "000011101100101001", xin_1 => "000011001101010001", pass => true),
  (xin_0 => "001001110100010001", xin_1 => "000111110001100111", pass => true),
  (xin_0 => "001011000001100101", xin_1 => "001010001100000001", pass => false),
  (xin_0 => "000111010000111100", xin_1 => "000011000001100011", pass => false),
  (xin_0 => "000111101011100001", xin_1 => "001010011001001011", pass => false),
  (xin_0 => "001001110100100110", xin_1 => "000010101001001101", pass => false),
  (xin_0 => "000110101100011110", xin_1 => "000011000100010001", pass => false),
  (xin_0 => "000110011011010111", xin_1 => "000100110100111100", pass => true),
  (xin_0 => "001010001000110001", xin_1 => "001010100111110010", pass => false),
  (xin_0 => "001000011011111011", xin_1 => "000010101110111000", pass => false),
  (xin_0 => "001001100011110001", xin_1 => "000100110101111110", pass => true),
  (xin_0 => "000101110111110011", xin_1 => "000010111111000001", pass => false),
  (xin_0 => "001001000011000110", xin_1 => "001001111011010110", pass => false),
  (xin_0 => "001100100101111110", xin_1 => "000111001001111110", pass => false),
  (xin_0 => "000110100111010011", xin_1 => "001001001111100001", pass => false),
  (xin_0 => "001100110011101010", xin_1 => "001010100010110010", pass => true),
  (xin_0 => "001101100110001011", xin_1 => "000110011000000010", pass => false),
  (xin_0 => "001111110101001110", xin_1 => "001001011111011001", pass => true),
  (xin_0 => "001011101010000110", xin_1 => "001001111001101011", pass => false),
  (xin_0 => "001011110101100000", xin_1 => "000111110000001010", pass => false),
  (xin_0 => "000101011010010111", xin_1 => "000110110000111110", pass => true),
  (xin_0 => "001011110010000000", xin_1 => "000001100101011110", pass => true),
  (xin_0 => "001010010111011001", xin_1 => "000101110101010110", pass => true),
  (xin_0 => "001100010111111001", xin_1 => "000110011110011111", pass => false),
  (xin_0 => "001011100011010110", xin_1 => "001000011111000000", pass => false),
  (xin_0 => "000110100010101101", xin_1 => "000010001100010000", pass => false),
  (xin_0 => "001100010001001010", xin_1 => "001000110111000011", pass => false),
  (xin_0 => "001100101111101000", xin_1 => "000000101111001000", pass => true),
  (xin_0 => "000110000110101001", xin_1 => "001001100101011111", pass => false),
  (xin_0 => "001000111100000011", xin_1 => "001011100010111101", pass => false),
  (xin_0 => "001010010110110100", xin_1 => "001001011001000001", pass => false),
  (xin_0 => "000111000110100000", xin_1 => "000011011000000110", pass => false),
  (xin_0 => "000111101101110010", xin_1 => "000100110000000111", pass => true),
  (xin_0 => "001000111010110001", xin_1 => "001010100010000100", pass => false),
  (xin_0 => "001110101111111100", xin_1 => "001011011011000000", pass => true),
  (xin_0 => "000100100011100111", xin_1 => "001001000110101000", pass => false),
  (xin_0 => "000101011101001101", xin_1 => "001001110101101111", pass => false),
  (xin_0 => "000111010101000100", xin_1 => "000001111101000010", pass => false),
  (xin_0 => "000101010110001101", xin_1 => "001001101011110100", pass => false),
  (xin_0 => "001001001100110011", xin_1 => "000011101000110000", pass => false),
  (xin_0 => "000110011101101111", xin_1 => "001000111010110011", pass => false),
  (xin_0 => "001011101110100001", xin_1 => "000100011111010000", pass => true),
  (xin_0 => "000111010001000011", xin_1 => "000100011100011000", pass => true),
  (xin_0 => "001001010100011001", xin_1 => "000011100110010100", pass => false),
  (xin_0 => "001010010001011101", xin_1 => "000011100101100001", pass => true),
  (xin_0 => "001001110010100100", xin_1 => "001001010010011000", pass => false),
  (xin_0 => "000100000011101011", xin_1 => "000010110000111101", pass => true),
  (xin_0 => "001100010110110100", xin_1 => "001010000110110001", pass => false),
  (xin_0 => "000101011101110101", xin_1 => "000111011100011101", pass => true),
  (xin_0 => "000111010100000011", xin_1 => "000010001011110101", pass => false),
  (xin_0 => "001100110011011010", xin_1 => "000011111000000001", pass => true),
  (xin_0 => "001011101000001101", xin_1 => "001001000100000010", pass => false),
  (xin_0 => "001001011010101000", xin_1 => "000100010110110000", pass => true),
  (xin_0 => "000101010010110100", xin_1 => "000100101010011100", pass => true),
  (xin_0 => "000110001010010010", xin_1 => "000110100011101000", pass => true),
  (xin_0 => "000111110110011000", xin_1 => "000011010100000100", pass => false),
  (xin_0 => "001011001110101111", xin_1 => "001000110101101001", pass => false),
  (xin_0 => "000111111100101111", xin_1 => "000111111110010001", pass => true),
  (xin_0 => "000111011011110001", xin_1 => "000011100111111010", pass => false),
  (xin_0 => "000110001110011101", xin_1 => "001001001100011100", pass => false),
  (xin_0 => "001011110111111000", xin_1 => "000111100101001111", pass => false),
  (xin_0 => "000111011110111001", xin_1 => "001011111110110101", pass => false),
  (xin_0 => "001011010111011101", xin_1 => "000110000011100101", pass => true),
  (xin_0 => "000110000100011111", xin_1 => "000010000000001010", pass => false),
  (xin_0 => "001000000111100001", xin_1 => "000111011001100001", pass => true),
  (xin_0 => "001000010111101111", xin_1 => "001000000010011111", pass => true),
  (xin_0 => "001010010000100011", xin_1 => "000110001100111100", pass => true),
  (xin_0 => "000111101100111101", xin_1 => "001001101011000011", pass => false),
  (xin_0 => "001001111101011100", xin_1 => "000111011111001010", pass => true),
  (xin_0 => "000110110001010110", xin_1 => "001001110100000000", pass => false),
  (xin_0 => "001101101100001010", xin_1 => "111111101010111001", pass => true),
  (xin_0 => "001100000101011100", xin_1 => "000111011000000000", pass => false),
  (xin_0 => "000111101001010100", xin_1 => "001011011001010001", pass => false),
  (xin_0 => "001101001101101110", xin_1 => "001010011101111000", pass => true),
  (xin_0 => "001000000111101110", xin_1 => "000010111110110100", pass => false),
  (xin_0 => "001000001000010101", xin_1 => "000011001000101001", pass => false),
  (xin_0 => "001010001000100110", xin_1 => "000110011011101010", pass => true),
  (xin_0 => "001100100111001110", xin_1 => "000110100000001001", pass => false),
  (xin_0 => "000101110111000000", xin_1 => "000100000100100110", pass => true),
  (xin_0 => "001000011011000010", xin_1 => "001001101101011011", pass => false),
  (xin_0 => "001010101100101110", xin_1 => "001001011101001110", pass => false),
  (xin_0 => "000110111011000110", xin_1 => "000010011011100000", pass => false),
  (xin_0 => "000100001101111001", xin_1 => "000111110100100010", pass => false),
  (xin_0 => "001110010001111100", xin_1 => "001001110011111110", pass => true),
  (xin_0 => "001001101100000101", xin_1 => "000011100110110101", pass => false),
  (xin_0 => "001100010001011101", xin_1 => "000110111101110001", pass => false),
  (xin_0 => "001100011110111110", xin_1 => "000101001000010000", pass => true),
  (xin_0 => "000110001101110110", xin_1 => "000100010010010010", pass => true),
  (xin_0 => "000111110100110000", xin_1 => "000011001001111101", pass => false),
  (xin_0 => "000111000101000000", xin_1 => "000010100001100000", pass => false),
  (xin_0 => "001000100011011110", xin_1 => "000111100001001010", pass => true),
  (xin_0 => "001100000011001001", xin_1 => "000110000110001001", pass => false),
  (xin_0 => "001011011001110000", xin_1 => "000110001111111101", pass => true),
  (xin_0 => "000110101110101000", xin_1 => "000011000101001000", pass => false),
  (xin_0 => "001000001011000100", xin_1 => "000001110000110111", pass => false),
  (xin_0 => "001010111010000110", xin_1 => "001000010000010001", pass => false),
  (xin_0 => "001010100101001110", xin_1 => "000110101111111110", pass => true),
  (xin_0 => "000111000011010110", xin_1 => "000101001101100110", pass => true),
  (xin_0 => "000110111101001010", xin_1 => "000001110011101100", pass => false),
  (xin_0 => "001000011100010100", xin_1 => "000101100110010100", pass => true),
  (xin_0 => "000111001100110001", xin_1 => "000001100111001001", pass => false),
  (xin_0 => "000111001101111001", xin_1 => "001010000001001001", pass => false),
  (xin_0 => "000111001001110111", xin_1 => "001001110001000111", pass => false),
  (xin_0 => "000110001100000110", xin_1 => "001000110011100110", pass => false),
  (xin_0 => "001100101100101110", xin_1 => "001000010010010111", pass => false),
  (xin_0 => "001000001000000101", xin_1 => "001010011100010000", pass => false),
  (xin_0 => "001101110100110111", xin_1 => "000101010000010000", pass => false),
  (xin_0 => "000110010000100010", xin_1 => "000100101100110101", pass => true),
  (xin_0 => "000100001100111010", xin_1 => "000010101100111101", pass => true),
  (xin_0 => "001100110110111011", xin_1 => "001010010000110111", pass => true),
  (xin_0 => "001011001011100111", xin_1 => "001000110100110101", pass => false),
  (xin_0 => "001000011100101001", xin_1 => "000011010110100111", pass => false),
  (xin_0 => "000100011000110111", xin_1 => "000111000011100011", pass => false),
  (xin_0 => "001000110110101110", xin_1 => "001010110110101101", pass => false),
  (xin_0 => "001010101111011101", xin_1 => "000100011100110001", pass => true),
  (xin_0 => "000100101101111101", xin_1 => "000110011110101100", pass => true),
  (xin_0 => "001001110010000110", xin_1 => "001001111101101000", pass => false),
  (xin_0 => "001000100111001101", xin_1 => "000010011001110100", pass => false),
  (xin_0 => "000111100011101010", xin_1 => "000100110000001010", pass => true),
  (xin_0 => "001010110111101010", xin_1 => "000110010001011011", pass => true),
  (xin_0 => "001010101101000001", xin_1 => "000100000100100011", pass => true),
  (xin_0 => "001010111011100101", xin_1 => "000110000111110100", pass => true),
  (xin_0 => "001000000010110010", xin_1 => "000011001111000011", pass => false),
  (xin_0 => "001101011011010100", xin_1 => "000101011011111100", pass => false),
  (xin_0 => "000100011111111010", xin_1 => "000100010001111100", pass => true),
  (xin_0 => "001001111010011101", xin_1 => "000110110010100000", pass => true),
  (xin_0 => "000111100000111110", xin_1 => "001001010110101101", pass => false),
  (xin_0 => "000100000000111001", xin_1 => "000100100010110111", pass => true),
  (xin_0 => "000110101100001101", xin_1 => "000101111000100010", pass => true),
  (xin_0 => "001010110111111110", xin_1 => "001011011000010110", pass => false),
  (xin_0 => "001000111110001111", xin_1 => "000110010000110111", pass => true),
  (xin_0 => "001011100100010101", xin_1 => "000010111100110100", pass => true),
  (xin_0 => "001000111010000011", xin_1 => "000100110111100000", pass => true),
  (xin_0 => "000110010010110000", xin_1 => "001001101011000001", pass => false),
  (xin_0 => "001000001001001111", xin_1 => "000101111100100001", pass => true),
  (xin_0 => "000110000110100110", xin_1 => "001001010110010101", pass => false),
  (xin_0 => "000111101100011101", xin_1 => "001101000010001110", pass => false),
  (xin_0 => "000111000110010100", xin_1 => "000101100000010100", pass => true),
  (xin_0 => "000101000100111111", xin_1 => "001000000010010010", pass => false),
  (xin_0 => "000100110111011101", xin_1 => "000011101000000100", pass => true),
  (xin_0 => "000110100010010010", xin_1 => "000010000110000100", pass => false),
  (xin_0 => "000111101100001010", xin_1 => "000011010101000010", pass => false),
  (xin_0 => "000110101010010010", xin_1 => "000010011010011010", pass => false),
  (xin_0 => "001011100110000011", xin_1 => "001100100110001100", pass => false),
  (xin_0 => "001011011101110001", xin_1 => "001000101100001000", pass => false),
  (xin_0 => "000110011001111000", xin_1 => "000010010110111101", pass => false),
  (xin_0 => "001001000111000111", xin_1 => "001100010100001101", pass => false),
  (xin_0 => "000111001001000100", xin_1 => "000100001011001100", pass => false),
  (xin_0 => "000111011010011001", xin_1 => "000110110001110101", pass => true),
  (xin_0 => "001000000101000011", xin_1 => "000010100001001010", pass => false),
  (xin_0 => "000100001000110101", xin_1 => "001000100000011001", pass => false),
  (xin_0 => "001010000001100011", xin_1 => "001001010111101011", pass => false),
  (xin_0 => "001010111110111000", xin_1 => "001001101100101000", pass => false),
  (xin_0 => "001010101111000100", xin_1 => "000111111011000010", pass => false),
  (xin_0 => "000110010101011100", xin_1 => "000101100111001010", pass => true),
  (xin_0 => "001011010101100000", xin_1 => "000111110000000001", pass => false),
  (xin_0 => "000101101001011101", xin_1 => "001000010101011001", pass => false),
  (xin_0 => "000100100100000101", xin_1 => "000110110111111101", pass => true),
  (xin_0 => "001011101100110000", xin_1 => "001001001110001101", pass => false),
  (xin_0 => "000101000101110010", xin_1 => "000011100111000100", pass => true),
  (xin_0 => "001010000000011101", xin_1 => "000101011010001001", pass => true),
  (xin_0 => "001001010011100000", xin_1 => "001011001011111000", pass => false),
  (xin_0 => "001010101001001110", xin_1 => "001000010010100101", pass => false),
  (xin_0 => "001001010111100101", xin_1 => "000111000001101000", pass => true),
  (xin_0 => "000101011010001011", xin_1 => "000110011110110100", pass => true),
  (xin_0 => "000111101111010000", xin_1 => "001010011111101101", pass => false),
  (xin_0 => "001000001011111000", xin_1 => "001010001000010111", pass => false),
  (xin_0 => "001010101110110100", xin_1 => "000100000101011010", pass => true),
  (xin_0 => "000011101101110011", xin_1 => "000100100100111001", pass => true),
  (xin_0 => "001010010111001110", xin_1 => "001001001111010101", pass => false),
  (xin_0 => "001101001101001010", xin_1 => "000101111110001111", pass => false),
  (xin_0 => "000110100000101010", xin_1 => "000010110000010101", pass => false),
  (xin_0 => "001011100111000100", xin_1 => "000110111011011110", pass => false),
  (xin_0 => "001000110001100111", xin_1 => "000111001000101010", pass => true),
  (xin_0 => "001101101010110011", xin_1 => "000100111010110111", pass => false),
  (xin_0 => "001011110111101110", xin_1 => "000011111101111101", pass => true),
  (xin_0 => "000011111000100000", xin_1 => "000111001100010111", pass => false),
  (xin_0 => "000111011000111110", xin_1 => "000111000111010011", pass => true),
  (xin_0 => "000110111001000100", xin_1 => "000010110010110100", pass => false),
  (xin_0 => "000101110001101110", xin_1 => "001001110000111001", pass => false),
  (xin_0 => "000011011110100110", xin_1 => "000010101100001001", pass => true),
  (xin_0 => "000111011001101001", xin_1 => "001001011010010111", pass => false),
  (xin_0 => "001100011001110010", xin_1 => "000001001001000110", pass => true),
  (xin_0 => "001101001001001011", xin_1 => "000101101001111010", pass => false),
  (xin_0 => "000110000001111011", xin_1 => "000111010011111100", pass => true),
  (xin_0 => "000111101110110010", xin_1 => "000101011111101110", pass => true),
  (xin_0 => "001011110001100100", xin_1 => "001000111101010000", pass => false),
  (xin_0 => "000101110011100101", xin_1 => "000111100011101001", pass => true),
  (xin_0 => "000110011110001110", xin_1 => "000101100000111010", pass => true),
  (xin_0 => "001010001000101111", xin_1 => "001001101111100000", pass => false),
  (xin_0 => "001010000111110011", xin_1 => "000011001100100101", pass => false),
  (xin_0 => "001000101001111010", xin_1 => "000100111101111100", pass => true),
  (xin_0 => "000110110001000010", xin_1 => "000010111001110010", pass => false),
  (xin_0 => "001101000001110010", xin_1 => "000010000010111001", pass => true),
  (xin_0 => "001000100010010100", xin_1 => "001011010101000011", pass => false),
  (xin_0 => "000110101001011101", xin_1 => "000001010001111101", pass => false),
  (xin_0 => "001111000111000010", xin_1 => "001001011111000011", pass => true),
  (xin_0 => "001100000011000101", xin_1 => "001010111000101101", pass => false),
  (xin_0 => "000111100111100010", xin_1 => "000010111101101100", pass => false),
  (xin_0 => "001010001011110010", xin_1 => "000010100011110100", pass => false),
  (xin_0 => "001001111100110110", xin_1 => "001000111111001000", pass => false),
  (xin_0 => "000101101000100001", xin_1 => "000111011101100001", pass => true),
  (xin_0 => "001100100110110010", xin_1 => "000001011101000011", pass => true),
  (xin_0 => "001110110101101001", xin_1 => "001001001101111011", pass => true),
  (xin_0 => "000110110100001010", xin_1 => "001001010011010111", pass => false),
  (xin_0 => "000110000001100111", xin_1 => "000101110000011001", pass => true),
  (xin_0 => "001100010111001000", xin_1 => "001000000110000100", pass => false),
  (xin_0 => "001100001011000110", xin_1 => "000110000010010110", pass => false),
  (xin_0 => "001010010111100011", xin_1 => "001010001110000011", pass => false),
  (xin_0 => "000111110110100000", xin_1 => "000010001010001000", pass => false),
  (xin_0 => "000111001000000001", xin_1 => "000011100101111100", pass => false),
  (xin_0 => "000010110110011011", xin_1 => "000001101001000011", pass => true),
  (xin_0 => "001010001000100001", xin_1 => "001011101100110010", pass => false),
  (xin_0 => "000101000000011011", xin_1 => "001001001100010110", pass => false),
  (xin_0 => "001010100101111101", xin_1 => "000011010000011101", pass => true),
  (xin_0 => "001101010100001101", xin_1 => "001010110111000110", pass => true),
  (xin_0 => "001100111110100010", xin_1 => "000010110111100010", pass => true),
  (xin_0 => "000110011110010111", xin_1 => "000010001100001000", pass => false),
  (xin_0 => "001010111110011001", xin_1 => "000100001111000111", pass => true),
  (xin_0 => "000101111010111001", xin_1 => "001001001010100010", pass => false),
  (xin_0 => "000111011101111110", xin_1 => "000011010100111001", pass => false),
  (xin_0 => "001100001000110111", xin_1 => "000101010001101000", pass => true),
  (xin_0 => "001000011010011000", xin_1 => "000101011010100111", pass => true),
  (xin_0 => "001001111010100100", xin_1 => "000100001000011000", pass => true),
  (xin_0 => "000111010011111010", xin_1 => "000001000100000010", pass => false),
  (xin_0 => "001100001000011000", xin_1 => "000110101000000110", pass => false),
  (xin_0 => "001001100110000101", xin_1 => "000110101011010000", pass => true),
  (xin_0 => "001010000011001101", xin_1 => "001010011000010011", pass => false),
  (xin_0 => "000111001110001000", xin_1 => "001001111011111110", pass => false),
  (xin_0 => "000111011011010011", xin_1 => "000010000010011001", pass => false),
  (xin_0 => "001011110111111110", xin_1 => "001000101111111000", pass => false),
  (xin_0 => "000110001100010011", xin_1 => "001001011100000101", pass => false),
  (xin_0 => "000111101000101011", xin_1 => "001000110111011110", pass => false),
  (xin_0 => "000100010110111100", xin_1 => "000111001101010011", pass => false),
  (xin_0 => "001011100100101101", xin_1 => "001001011000011010", pass => false),
  (xin_0 => "000101101011010001", xin_1 => "000110101110011001", pass => true),
  (xin_0 => "000110011010101000", xin_1 => "000011001011100010", pass => false),
  (xin_0 => "000101011101011100", xin_1 => "000101000010001111", pass => true),
  (xin_0 => "001010011001110110", xin_1 => "000110010011011101", pass => true),
  (xin_0 => "000110010001000011", xin_1 => "000100011010101110", pass => true),
  (xin_0 => "000101101001110101", xin_1 => "000011011010010000", pass => true),
  (xin_0 => "001010000100110001", xin_1 => "000110001110011100", pass => true),
  (xin_0 => "001100000010011111", xin_1 => "000111100100101101", pass => false),
  (xin_0 => "001010101101001100", xin_1 => "001010000110110100", pass => false),
  (xin_0 => "001011010010010100", xin_1 => "000111100000001110", pass => false),
  (xin_0 => "001101101100010000", xin_1 => "001001100111100000", pass => true),
  (xin_0 => "001010001111110100", xin_1 => "000010101001001001", pass => false),
  (xin_0 => "000101101110000001", xin_1 => "000010101010001001", pass => false),
  (xin_0 => "000111100111111110", xin_1 => "000010110110001100", pass => false),
  (xin_0 => "001111101111101011", xin_1 => "001001110100000011", pass => true),
  (xin_0 => "001110011011010101", xin_1 => "001001100100001101", pass => true),
  (xin_0 => "000100000111101001", xin_1 => "000001101011000101", pass => true),
  (xin_0 => "001101111010111100", xin_1 => "001001100100110010", pass => true),
  (xin_0 => "001000010101011101", xin_1 => "001000100100011001", pass => true),
  (xin_0 => "000011010110011100", xin_1 => "001001001001010000", pass => false),
  (xin_0 => "000011110011001110", xin_1 => "000001011010011011", pass => true),
  (xin_0 => "000101010000101001", xin_1 => "000110110010010011", pass => true),
  (xin_0 => "000011110111110001", xin_1 => "000001010001111001", pass => true),
  (xin_0 => "001001110100110000", xin_1 => "001100010110001110", pass => false),
  (xin_0 => "000111101000001101", xin_1 => "000011001111011010", pass => false),
  (xin_0 => "000101101000000010", xin_1 => "001000011100010110", pass => false),
  (xin_0 => "001010010111010100", xin_1 => "001010101001011011", pass => false),
  (xin_0 => "001001011011011010", xin_1 => "000010101001010101", pass => false),
  (xin_0 => "001000100110011111", xin_1 => "000100101101101101", pass => true),
  (xin_0 => "000111010100100101", xin_1 => "000101101110101110", pass => true),
  (xin_0 => "000100100010110000", xin_1 => "001001000100001011", pass => false),
  (xin_0 => "000011100010000010", xin_1 => "000100110110110000", pass => true),
  (xin_0 => "001011101111001001", xin_1 => "000111100110111101", pass => false),
  (xin_0 => "000011110111100001", xin_1 => "000011011110110100", pass => true),
  (xin_0 => "001101000100111011", xin_1 => "000111010111010010", pass => false),
  (xin_0 => "001100011111010010", xin_1 => "000101111010000001", pass => false),
  (xin_0 => "001111000110101111", xin_1 => "001001001100110011", pass => true),
  (xin_0 => "001111010101010000", xin_1 => "000100001101001100", pass => false),
  (xin_0 => "000100100011011100", xin_1 => "000111110000111010", pass => false),
  (xin_0 => "000101001111011101", xin_1 => "000100100101000011", pass => true),
  (xin_0 => "001011000001010001", xin_1 => "001001000111000010", pass => false),
  (xin_0 => "000100010001000001", xin_1 => "000000100110101110", pass => true),
  (xin_0 => "001001010011011100", xin_1 => "000010010001101100", pass => false),
  (xin_0 => "000110101110111011", xin_1 => "001001011100110011", pass => false),
  (xin_0 => "001000110000110110", xin_1 => "001010000000001111", pass => false),
  (xin_0 => "001100000100110111", xin_1 => "001000011010101110", pass => false),
  (xin_0 => "001001010100101000", xin_1 => "001001111011110010", pass => false),
  (xin_0 => "001100010001010011", xin_1 => "000110110111110101", pass => false),
  (xin_0 => "000101110001100100", xin_1 => "001000101100010101", pass => false),
  (xin_0 => "001000001011011100", xin_1 => "000011100000001010", pass => false),
  (xin_0 => "001010101110101000", xin_1 => "000110000001111010", pass => true),
  (xin_0 => "001000101011101110", xin_1 => "000111101010011110", pass => true),
  (xin_0 => "001001101010111000", xin_1 => "000101100001010001", pass => true),
  (xin_0 => "001011110111001011", xin_1 => "001001110010110001", pass => false),
  (xin_0 => "000111000010111110", xin_1 => "000010010000010101", pass => false),
  (xin_0 => "001100010110000010", xin_1 => "000111100001100001", pass => false),
  (xin_0 => "001010011101011000", xin_1 => "001001111001110111", pass => false),
  (xin_0 => "001100000001010011", xin_1 => "001001000000010000", pass => false),
  (xin_0 => "001001100001010101", xin_1 => "001010000101101010", pass => false),
  (xin_0 => "001000011111101111", xin_1 => "000010111011101111", pass => false),
  (xin_0 => "001100101101101010", xin_1 => "001000001100101001", pass => false),
  (xin_0 => "001001101110001000", xin_1 => "000101000101100111", pass => true),
  (xin_0 => "000100000100010011", xin_1 => "000000100010011000", pass => true),
  (xin_0 => "001011000101010011", xin_1 => "000111111101100101", pass => false),
  (xin_0 => "000111110011011000", xin_1 => "000111111100000111", pass => true),
  (xin_0 => "001100011111110110", xin_1 => "000111111011110001", pass => false),
  (xin_0 => "001001100101111001", xin_1 => "000010000110011001", pass => false),
  (xin_0 => "000101001111110001", xin_1 => "000010101011101001", pass => true),
  (xin_0 => "001000100100011111", xin_1 => "000010000111011001", pass => false),
  (xin_0 => "001011001101010111", xin_1 => "000100000111011111", pass => true),
  (xin_0 => "001010001001011110", xin_1 => "000101110110100000", pass => true),
  (xin_0 => "000111010001101001", xin_1 => "000101000001010101", pass => true),
  (xin_0 => "000111001011101001", xin_1 => "000010010110000101", pass => false),
  (xin_0 => "001001011101111010", xin_1 => "000010000011011100", pass => false),
  (xin_0 => "001000010100000011", xin_1 => "000110100101111111", pass => true),
  (xin_0 => "000110111011110001", xin_1 => "000001000101101110", pass => false),
  (xin_0 => "001110011010111000", xin_1 => "000100010011011000", pass => false),
  (xin_0 => "000111100100000110", xin_1 => "001000111111101010", pass => false),
  (xin_0 => "000011100001011101", xin_1 => "000010111000110010", pass => true),
  (xin_0 => "001011010001110100", xin_1 => "000110101000011000", pass => false),
  (xin_0 => "001100100011001110", xin_1 => "000010001011110001", pass => true),
  (xin_0 => "000110000111101000", xin_1 => "001001000011101011", pass => false),
  (xin_0 => "001011010011011000", xin_1 => "001100010011110101", pass => false),
  (xin_0 => "000101001010001101", xin_1 => "001010000000111011", pass => false),
  (xin_0 => "000100001110010100", xin_1 => "001000011100001010", pass => false),
  (xin_0 => "001001011110111110", xin_1 => "000010100011001101", pass => false),
  (xin_0 => "001101011010001000", xin_1 => "000101101000111011", pass => false),
  (xin_0 => "000100000001000011", xin_1 => "001000110111100110", pass => false),
  (xin_0 => "001000010010010010", xin_1 => "001001100000111110", pass => false),
  (xin_0 => "001011001000010000", xin_1 => "001000000100110111", pass => false),
  (xin_0 => "000100110100100001", xin_1 => "001010000100000001", pass => false),
  (xin_0 => "001010001101011110", xin_1 => "000101101001110010", pass => true),
  (xin_0 => "001000100001011101", xin_1 => "000110001010111110", pass => true),
  (xin_0 => "001100000110000101", xin_1 => "000110001110011010", pass => false),
  (xin_0 => "001101111000100001", xin_1 => "000110101101001000", pass => false),
  (xin_0 => "001001001001000000", xin_1 => "000010100001111000", pass => false),
  (xin_0 => "000100110111001011", xin_1 => "001001100110010001", pass => false),
  (xin_0 => "001011110010010101", xin_1 => "000010001100010010", pass => true),
  (xin_0 => "000111101100100000", xin_1 => "000010111000000010", pass => false),
  (xin_0 => "001000111110101011", xin_1 => "000100111010001010", pass => true),
  (xin_0 => "001001111011001101", xin_1 => "000100110000100010", pass => true),
  (xin_0 => "001100100001011101", xin_1 => "000011110101110111", pass => true),
  (xin_0 => "000110111111101000", xin_1 => "001000101001100011", pass => false),
  (xin_0 => "001100010000010010", xin_1 => "000101100101111101", pass => true),
  (xin_0 => "001000101000111111", xin_1 => "001011011001100001", pass => false),
  (xin_0 => "001000110100100101", xin_1 => "001011100010010111", pass => false),
  (xin_0 => "001011000110100001", xin_1 => "001000011111001110", pass => false),
  (xin_0 => "001000101100010111", xin_1 => "000101111000000110", pass => true),
  (xin_0 => "001011001000011000", xin_1 => "001011000001010011", pass => false),
  (xin_0 => "001100011110100111", xin_1 => "001001101010011111", pass => false),
  (xin_0 => "000111100000001010", xin_1 => "000110011101110111", pass => true),
  (xin_0 => "001000101111110111", xin_1 => "000111100011111001", pass => true),
  (xin_0 => "001011000100010110", xin_1 => "000011001101111000", pass => true),
  (xin_0 => "001100110110001111", xin_1 => "000101011011101110", pass => false),
  (xin_0 => "001100010000100000", xin_1 => "000111101110100101", pass => false),
  (xin_0 => "000100001001100100", xin_1 => "000011111111101000", pass => true),
  (xin_0 => "000101111111011010", xin_1 => "000010010100011011", pass => false),
  (xin_0 => "001100111100010010", xin_1 => "001000000000000000", pass => false),
  (xin_0 => "000110011001110000", xin_1 => "000111011101101011", pass => true),
  (xin_0 => "001000100111011111", xin_1 => "000110011110011010", pass => true),
  (xin_0 => "000111000000010100", xin_1 => "000110000110100000", pass => true),
  (xin_0 => "001010011001001001", xin_1 => "000100001100000000", pass => true),
  (xin_0 => "000110111010010000", xin_1 => "000011011001101010", pass => false),
  (xin_0 => "001001000111001110", xin_1 => "001010010100001100", pass => false),
  (xin_0 => "001000100000010101", xin_1 => "001010001010001000", pass => false),
  (xin_0 => "000110100001001010", xin_1 => "000011000011001111", pass => false),
  (xin_0 => "001001110011000010", xin_1 => "000011110011111001", pass => false),
  (xin_0 => "001011100011011000", xin_1 => "001001011110111110", pass => false),
  (xin_0 => "001010101001101101", xin_1 => "000111011100110111", pass => false),
  (xin_0 => "000101010101000010", xin_1 => "000001101111110011", pass => false),
  (xin_0 => "001001011000110110", xin_1 => "000111100100011101", pass => true),
  (xin_0 => "000110011001011001", xin_1 => "000100011000010101", pass => true),
  (xin_0 => "001010111011111111", xin_1 => "000111111000101101", pass => false),
  (xin_0 => "001010000010010101", xin_1 => "001001001010100001", pass => false),
  (xin_0 => "001100111111100011", xin_1 => "000111110000101100", pass => false),
  (xin_0 => "001100101111110110", xin_1 => "000101100000001111", pass => false),
  (xin_0 => "001001100100110110", xin_1 => "000001001011110011", pass => false),
  (xin_0 => "001001101111100011", xin_1 => "001011101010100101", pass => false),
  (xin_0 => "001001101110110110", xin_1 => "001000000100010100", pass => true),
  (xin_0 => "001010011001001000", xin_1 => "001101000000000010", pass => false),
  (xin_0 => "001011111110011110", xin_1 => "000111000101111101", pass => false),
  (xin_0 => "001001100101000010", xin_1 => "000010110011110101", pass => false),
  (xin_0 => "000100010000110000", xin_1 => "000011100000010110", pass => true),
  (xin_0 => "010000011111101101", xin_1 => "001001000111100010", pass => true),
  (xin_0 => "000101001110111110", xin_1 => "000110001101100110", pass => true),
  (xin_0 => "001000011100010001", xin_1 => "001010110100000101", pass => false),
  (xin_0 => "001011001110100110", xin_1 => "000110110000001110", pass => false),
  (xin_0 => "001010011100110100", xin_1 => "001010101011000011", pass => false),
  (xin_0 => "001010111010100000", xin_1 => "001001010110101100", pass => false),
  (xin_0 => "001100000100010010", xin_1 => "000111100100010110", pass => false),
  (xin_0 => "001010010110111101", xin_1 => "001000001010000110", pass => false),
  (xin_0 => "001000011111111001", xin_1 => "001011110101001000", pass => false),
  (xin_0 => "000111010010001000", xin_1 => "000100110100100011", pass => true),
  (xin_0 => "000100100001101100", xin_1 => "000010101011101100", pass => true),
  (xin_0 => "001101100001100001", xin_1 => "000110110110101101", pass => false),
  (xin_0 => "001001101110000100", xin_1 => "000101101011000101", pass => true),
  (xin_0 => "000100000011000110", xin_1 => "000010100101110011", pass => true),
  (xin_0 => "000111011000011011", xin_1 => "000011111110101110", pass => false),
  (xin_0 => "000110101101111000", xin_1 => "000010000010011010", pass => false),
  (xin_0 => "001000001101000000", xin_1 => "001001010000011000", pass => false),
  (xin_0 => "000111101001011001", xin_1 => "000010001010101110", pass => false),
  (xin_0 => "001001111000011111", xin_1 => "001011000010110001", pass => false),
  (xin_0 => "000101000100111000", xin_1 => "001000011010000001", pass => false),
  (xin_0 => "000100011001111100", xin_1 => "000001110000101001", pass => true),
  (xin_0 => "001010010000100110", xin_1 => "000010011110010011", pass => false),
  (xin_0 => "001011010001010100", xin_1 => "001000001111010000", pass => false),
  (xin_0 => "001001011110000010", xin_1 => "001010110000100111", pass => false),
  (xin_0 => "000011100100010110", xin_1 => "000010010001001100", pass => true),
  (xin_0 => "001001000010100110", xin_1 => "000011100000100011", pass => false),
  (xin_0 => "000100100101000000", xin_1 => "000111101100001110", pass => false),
  (xin_0 => "001000100111011010", xin_1 => "000010011110111111", pass => false),
  (xin_0 => "000101110011111010", xin_1 => "000011100101101110", pass => true),
  (xin_0 => "001001011010001001", xin_1 => "001001001000100101", pass => false),
  (xin_0 => "000100111000111001", xin_1 => "001001001101001000", pass => false),
  (xin_0 => "000010110100000010", xin_1 => "000100011110101101", pass => true),
  (xin_0 => "000110101100100101", xin_1 => "001001100010011001", pass => false),
  (xin_0 => "001001011011110000", xin_1 => "000101001110011000", pass => true),
  (xin_0 => "001011011101100110", xin_1 => "000011110001100100", pass => true),
  (xin_0 => "001011011010100111", xin_1 => "000011101101010010", pass => true),
  (xin_0 => "001001100110111001", xin_1 => "000011001000011001", pass => false),
  (xin_0 => "001001011011001100", xin_1 => "000010111101000010", pass => false),
  (xin_0 => "000111101111110010", xin_1 => "000011010111011110", pass => false),
  (xin_0 => "000100110111010011", xin_1 => "000101100100111010", pass => true),
  (xin_0 => "001101100011100110", xin_1 => "000101000101000010", pass => false),
  (xin_0 => "001010110101111001", xin_1 => "000100010000110111", pass => true),
  (xin_0 => "010000001111000110", xin_1 => "001000111101110100", pass => true),
  (xin_0 => "001000110111111010", xin_1 => "000001111011010000", pass => false),
  (xin_0 => "001101010111010111", xin_1 => "001000101001001001", pass => false),
  (xin_0 => "001000100110000101", xin_1 => "000010110100001001", pass => false),
  (xin_0 => "001100100100010110", xin_1 => "000010011010110000", pass => true),
  (xin_0 => "001001001010011001", xin_1 => "001011101101010011", pass => false),
  (xin_0 => "000111110111111110", xin_1 => "000010110111000111", pass => false),
  (xin_0 => "001001010110011111", xin_1 => "000101011110100101", pass => true),
  (xin_0 => "001000111101111110", xin_1 => "000110111101001111", pass => true),
  (xin_0 => "001011110000000101", xin_1 => "000101100111111010", pass => true),
  (xin_0 => "001010100011100010", xin_1 => "000101101111100100", pass => true),
  (xin_0 => "001000000110011000", xin_1 => "000111111100100100", pass => true),
  (xin_0 => "000111100000010111", xin_1 => "000110000010111110", pass => true),
  (xin_0 => "001001100001001001", xin_1 => "000101010101000000", pass => true),
  (xin_0 => "001100001011111101", xin_1 => "000100001110010100", pass => true),
  (xin_0 => "001000110000000101", xin_1 => "001010111101001111", pass => false),
  (xin_0 => "001000010011110000", xin_1 => "001101101110001100", pass => false),
  (xin_0 => "001100101100001111", xin_1 => "000110010111000100", pass => false),
  (xin_0 => "001000010011110010", xin_1 => "000111000000111110", pass => true),
  (xin_0 => "000110110111101011", xin_1 => "000110111101101010", pass => true),
  (xin_0 => "001000101001001001", xin_1 => "000101100001011000", pass => true),
  (xin_0 => "000110011010101111", xin_1 => "001000000001100101", pass => true),
  (xin_0 => "001000001100111001", xin_1 => "001010110110110111", pass => false),
  (xin_0 => "001011010011110010", xin_1 => "001001011101011111", pass => false),
  (xin_0 => "000011101111101111", xin_1 => "000001000001111000", pass => true),
  (xin_0 => "001010011000101010", xin_1 => "001001110011001011", pass => false),
  (xin_0 => "001100010111101110", xin_1 => "001000000000011000", pass => false),
  (xin_0 => "000101101011111100", xin_1 => "000110000010001110", pass => true),
  (xin_0 => "000111011111100110", xin_1 => "001001010110001010", pass => false),
  (xin_0 => "001000110011100011", xin_1 => "000011010001011101", pass => false),
  (xin_0 => "001100110010111000", xin_1 => "001011011001001111", pass => true),
  (xin_0 => "001110000110000000", xin_1 => "000110111101001001", pass => false),
  (xin_0 => "001000011011110100", xin_1 => "000110000101000000", pass => true),
  (xin_0 => "000100100001100111", xin_1 => "000110010011011100", pass => true),
  (xin_0 => "001001001010011110", xin_1 => "000001110010000011", pass => false),
  (xin_0 => "001100000100111011", xin_1 => "000111100011011111", pass => false),
  (xin_0 => "000111111101101001", xin_1 => "000010001111010110", pass => false),
  (xin_0 => "001010010110000000", xin_1 => "000010111000000101", pass => false),
  (xin_0 => "000100001110100011", xin_1 => "000010101101101010", pass => true),
  (xin_0 => "010000100101101100", xin_1 => "001001001010011011", pass => true),
  (xin_0 => "001001010010110101", xin_1 => "000010000100010111", pass => false),
  (xin_0 => "001011010111101101", xin_1 => "000100011101000000", pass => true),
  (xin_0 => "001100001110111010", xin_1 => "000111011101010011", pass => false),
  (xin_0 => "000101010100111110", xin_1 => "000010010110000011", pass => false),
  (xin_0 => "001100010000011100", xin_1 => "001000101100111011", pass => false),
  (xin_0 => "001100100011001000", xin_1 => "000111000011101101", pass => false),
  (xin_0 => "001010000101011101", xin_1 => "000001111011000011", pass => false),
  (xin_0 => "000011010100110110", xin_1 => "000011111010011110", pass => true),
  (xin_0 => "001010110011110001", xin_1 => "001010010101100111", pass => false),
  (xin_0 => "000100101111110000", xin_1 => "000101101110000110", pass => true),
  (xin_0 => "001010100000101110", xin_1 => "000010011010101101", pass => false),
  (xin_0 => "000111001100001000", xin_1 => "000011011100010000", pass => false),
  (xin_0 => "001001110100001111", xin_1 => "000011100011110011", pass => false),
  (xin_0 => "000100100000010100", xin_1 => "000111111011111101", pass => false),
  (xin_0 => "001101101100110011", xin_1 => "001010101011000111", pass => true),
  (xin_0 => "000111011010001011", xin_1 => "000101000000010100", pass => true),
  (xin_0 => "001011010011011100", xin_1 => "000001001110000001", pass => true),
  (xin_0 => "000111110010010001", xin_1 => "000100101111100111", pass => true),
  (xin_0 => "001011100100101101", xin_1 => "001001101110101111", pass => false),
  (xin_0 => "001101010000100101", xin_1 => "001000001000100100", pass => false),
  (xin_0 => "000111110010110101", xin_1 => "000110001111011101", pass => true),
  (xin_0 => "000101111001000000", xin_1 => "001001010111001001", pass => false),
  (xin_0 => "001011011000100110", xin_1 => "000101111110101000", pass => true),
  (xin_0 => "000101010001010000", xin_1 => "000100001011100010", pass => true),
  (xin_0 => "000110011101010110", xin_1 => "000011100110110100", pass => false),
  (xin_0 => "000111011101100000", xin_1 => "001001001100011100", pass => false),
  (xin_0 => "001000110000110010", xin_1 => "000010001011111011", pass => false),
  (xin_0 => "001011111010101011", xin_1 => "001000110101011010", pass => false),
  (xin_0 => "001011011110111001", xin_1 => "000011000110011011", pass => true),
  (xin_0 => "001010010001110111", xin_1 => "000100000100101000", pass => true),
  (xin_0 => "001000101010010100", xin_1 => "000101110110111010", pass => true),
  (xin_0 => "001000101100000111", xin_1 => "000101111110001001", pass => true),
  (xin_0 => "000101000011010101", xin_1 => "000010100110011101", pass => true),
  (xin_0 => "001000001011110000", xin_1 => "000010100101100011", pass => false),
  (xin_0 => "001000111111010111", xin_1 => "001010001010000001", pass => false),
  (xin_0 => "001011100010101101", xin_1 => "000011111110001010", pass => true),
  (xin_0 => "001000011111000010", xin_1 => "000110001010001110", pass => true),
  (xin_0 => "000100100001010000", xin_1 => "000010100011100010", pass => true),
  (xin_0 => "001000111010010111", xin_1 => "001010111011001011", pass => false),
  (xin_0 => "000110100010000010", xin_1 => "000100101011111101", pass => true),
  (xin_0 => "001000111001011101", xin_1 => "000011000101100101", pass => false),
  (xin_0 => "001000111110100111", xin_1 => "000011011100000011", pass => false),
  (xin_0 => "000111100011110011", xin_1 => "001001100010010111", pass => false),
  (xin_0 => "010000000001001111", xin_1 => "000100110111011010", pass => false),
  (xin_0 => "001000000101101010", xin_1 => "000101011111011000", pass => true),
  (xin_0 => "001100111011001111", xin_1 => "001010001010010110", pass => true),
  (xin_0 => "001010001001100011", xin_1 => "000010010001010111", pass => false),
  (xin_0 => "001001001101010011", xin_1 => "000010111100010011", pass => false),
  (xin_0 => "001010111001111010", xin_1 => "001101111000010000", pass => false),
  (xin_0 => "000100000111100011", xin_1 => "000110001101101100", pass => true),
  (xin_0 => "001010100110111110", xin_1 => "000001100101101110", pass => false),
  (xin_0 => "001001010101001100", xin_1 => "001010011011100100", pass => false),
  (xin_0 => "001011010100010101", xin_1 => "001000100010101110", pass => false),
  (xin_0 => "001101100000010110", xin_1 => "001010100101101101", pass => true),
  (xin_0 => "001000111110101101", xin_1 => "000111100010011101", pass => true),
  (xin_0 => "001011000100000000", xin_1 => "001000100000110111", pass => false),
  (xin_0 => "001001000010011011", xin_1 => "000010100010100101", pass => false),
  (xin_0 => "001010000100111100", xin_1 => "001000110110100000", pass => false),
  (xin_0 => "001011010011100000", xin_1 => "000011111100100010", pass => true),
  (xin_0 => "001001100100011111", xin_1 => "000011111100010011", pass => false),
  (xin_0 => "000100010010101000", xin_1 => "000101000111110001", pass => true),
  (xin_0 => "001000111001010100", xin_1 => "000010001110001000", pass => false),
  (xin_0 => "000110101011100000", xin_1 => "000010110101101100", pass => false),
  (xin_0 => "000110000010011000", xin_1 => "001001111010110011", pass => false),
  (xin_0 => "001011010001001101", xin_1 => "000011101100010001", pass => true),
  (xin_0 => "001010011101101011", xin_1 => "000111010111100110", pass => true),
  (xin_0 => "001000110000111010", xin_1 => "001000001001001110", pass => true),
  (xin_0 => "001100100100101000", xin_1 => "000010000010110101", pass => true),
  (xin_0 => "001010000110010001", xin_1 => "001001111001001100", pass => false),
  (xin_0 => "010000001101101011", xin_1 => "001010001011011011", pass => true),
  (xin_0 => "001011010101100101", xin_1 => "001001011000100011", pass => false),
  (xin_0 => "001001101000100100", xin_1 => "000011000010011110", pass => false),
  (xin_0 => "000101110100000100", xin_1 => "000110100100101010", pass => true),
  (xin_0 => "001010100110011110", xin_1 => "001010100111010011", pass => false),
  (xin_0 => "001010011110101011", xin_1 => "000101011101101101", pass => true),
  (xin_0 => "000101110001111101", xin_1 => "001010011101101011", pass => false),
  (xin_0 => "000101110111001101", xin_1 => "000100110101110011", pass => true),
  (xin_0 => "001000110000100001", xin_1 => "001011110110110101", pass => false),
  (xin_0 => "001100100110111100", xin_1 => "000010000011001110", pass => true),
  (xin_0 => "001000101000101011", xin_1 => "000101000110010001", pass => true),
  (xin_0 => "000110101011101100", xin_1 => "000110001101010011", pass => true),
  (xin_0 => "001101100000101101", xin_1 => "000101111111010001", pass => false),
  (xin_0 => "001001010100110101", xin_1 => "000011100001101100", pass => false),
  (xin_0 => "001000111000001001", xin_1 => "000010101001010011", pass => false),
  (xin_0 => "000110010011111010", xin_1 => "001010010011010110", pass => false),
  (xin_0 => "001011011011011110", xin_1 => "000011101101101101", pass => true),
  (xin_0 => "000101100000111101", xin_1 => "000100010010011101", pass => true),
  (xin_0 => "000111010111100001", xin_1 => "001011011010011000", pass => false),
  (xin_0 => "000101011000010000", xin_1 => "000100000101110111", pass => true),
  (xin_0 => "000110001110010110", xin_1 => "000010101110011110", pass => false),
  (xin_0 => "001000001101000110", xin_1 => "000011000000101100", pass => false),
  (xin_0 => "000101110110000101", xin_1 => "000111110110010111", pass => true),
  (xin_0 => "001000010011100101", xin_1 => "001001011001000011", pass => false),
  (xin_0 => "001001000000101101", xin_1 => "000001100010010100", pass => false),
  (xin_0 => "000101111111001010", xin_1 => "001000010001111101", pass => false),
  (xin_0 => "000101001001000110", xin_1 => "001001010000000110", pass => false),
  (xin_0 => "000111001010100011", xin_1 => "000100110101011100", pass => true),
  (xin_0 => "000111100010101000", xin_1 => "000010100110001111", pass => false),
  (xin_0 => "001010011101111110", xin_1 => "001001011011010100", pass => false),
  (xin_0 => "000100000110000100", xin_1 => "000100110010101001", pass => true),
  (xin_0 => "001000011000010100", xin_1 => "000100100110010010", pass => true),
  (xin_0 => "001011000010100111", xin_1 => "000101110000101010", pass => true),
  (xin_0 => "001000011011111111", xin_1 => "000101100000001110", pass => true),
  (xin_0 => "001010000011001111", xin_1 => "001010010111100010", pass => false),
  (xin_0 => "001110000110001111", xin_1 => "001001110101110010", pass => true),
  (xin_0 => "000111100101111000", xin_1 => "000010110100011011", pass => false),
  (xin_0 => "001101001101110011", xin_1 => "000111101101001010", pass => false),
  (xin_0 => "001010110010011101", xin_1 => "001000111101111100", pass => false),
  (xin_0 => "001100000100010111", xin_1 => "000011001110110101", pass => true),
  (xin_0 => "001000000101100100", xin_1 => "000010110001000011", pass => false),
  (xin_0 => "001000110000011101", xin_1 => "000101000001111100", pass => true),
  (xin_0 => "000110101010100000", xin_1 => "000011101110100001", pass => false),
  (xin_0 => "000110111001111001", xin_1 => "000100100000000101", pass => true),
  (xin_0 => "001101001001000100", xin_1 => "000011000101010101", pass => true),
  (xin_0 => "001100101001111001", xin_1 => "000101001100010100", pass => true),
  (xin_0 => "000111110100011110", xin_1 => "001010001111010101", pass => false),
  (xin_0 => "001011010111101100", xin_1 => "000101101100001011", pass => true),
  (xin_0 => "000011111010111111", xin_1 => "001001001100001010", pass => false),
  (xin_0 => "001010001101001111", xin_1 => "000111011000100011", pass => true),
  (xin_0 => "000110001000101101", xin_1 => "000111101010100111", pass => true),
  (xin_0 => "001011011100001000", xin_1 => "000111011100001110", pass => false),
  (xin_0 => "001000110100000110", xin_1 => "000010111111100101", pass => false),
  (xin_0 => "001011101000001000", xin_1 => "000110111110010101", pass => false),
  (xin_0 => "001000011001110011", xin_1 => "000001111011000011", pass => false),
  (xin_0 => "000100111001011001", xin_1 => "000101000110100000", pass => true),
  (xin_0 => "000111110011111001", xin_1 => "000101001100110111", pass => true),
  (xin_0 => "001001010101110001", xin_1 => "000011000000100011", pass => false),
  (xin_0 => "000011001110011011", xin_1 => "000011100011011001", pass => true),
  (xin_0 => "001100110010100111", xin_1 => "000101110010100010", pass => false),
  (xin_0 => "001110001111001100", xin_1 => "001010100100110111", pass => true),
  (xin_0 => "000101110101001111", xin_1 => "000010000000101010", pass => false),
  (xin_0 => "001000110111011111", xin_1 => "000001011010110111", pass => false),
  (xin_0 => "001000100011011010", xin_1 => "000011010101101001", pass => false),
  (xin_0 => "000011010111110101", xin_1 => "000101010001010101", pass => true),
  (xin_0 => "001000010111011010", xin_1 => "001010000011011110", pass => false),
  (xin_0 => "001001111111010000", xin_1 => "000010111101110101", pass => false),
  (xin_0 => "000100011001000000", xin_1 => "000111011000000100", pass => false),
  (xin_0 => "000110010111110100", xin_1 => "001001010001000110", pass => false),
  (xin_0 => "000110110011111010", xin_1 => "001010010000010000", pass => false),
  (xin_0 => "000100111100010011", xin_1 => "000101110001101001", pass => true),
  (xin_0 => "000100001101010100", xin_1 => "000000011010101011", pass => true),
  (xin_0 => "001101011100110100", xin_1 => "000110001101100000", pass => false),
  (xin_0 => "001001110000110000", xin_1 => "000110101011100111", pass => true),
  (xin_0 => "001101101011110001", xin_1 => "000111101011000100", pass => false),
  (xin_0 => "001001111011000101", xin_1 => "001100001010101110", pass => false),
  (xin_0 => "000111100100000010", xin_1 => "000011011100111100", pass => false),
  (xin_0 => "001100101011010100", xin_1 => "000111010000001010", pass => false),
  (xin_0 => "001100101011011000", xin_1 => "000110101100000011", pass => false),
  (xin_0 => "001000101000111111", xin_1 => "000010010001010000", pass => false),
  (xin_0 => "001000100000101101", xin_1 => "000010101111100101", pass => false),
  (xin_0 => "000110111110011001", xin_1 => "001010011010010011", pass => false),
  (xin_0 => "001100001110100110", xin_1 => "001010101110011100", pass => false),
  (xin_0 => "000111000011111001", xin_1 => "000111100010110001", pass => true),
  (xin_0 => "000101101111110101", xin_1 => "000011101110110010", pass => true),
  (xin_0 => "000100100101111111", xin_1 => "000011101101010111", pass => true),
  (xin_0 => "001000101110100100", xin_1 => "000011010010011001", pass => false),
  (xin_0 => "001100000110111001", xin_1 => "000010110101001000", pass => true),
  (xin_0 => "001100011100000101", xin_1 => "001010111010010011", pass => true),
  (xin_0 => "001100110110101111", xin_1 => "000110111011001000", pass => false),
  (xin_0 => "000011010001001101", xin_1 => "000011010111010111", pass => true),
  (xin_0 => "001000010001111011", xin_1 => "000001111110110111", pass => false),
  (xin_0 => "000100011101011000", xin_1 => "000001011000010000", pass => true),
  (xin_0 => "000101100111011101", xin_1 => "001000100100100010", pass => false),
  (xin_0 => "001000000010011001", xin_1 => "000110110001000011", pass => true),
  (xin_0 => "001011000010010110", xin_1 => "000110011101110000", pass => true),
  (xin_0 => "001101100010110110", xin_1 => "000010010011101111", pass => true),
  (xin_0 => "001100110000010110", xin_1 => "000110101100000001", pass => false),
  (xin_0 => "001110001011011011", xin_1 => "001010010111011010", pass => true),
  (xin_0 => "000111001001011111", xin_1 => "001001111111110010", pass => false),
  (xin_0 => "001100110100110000", xin_1 => "000111000011111001", pass => false),
  (xin_0 => "001100000100010110", xin_1 => "000111100011110000", pass => false),
  (xin_0 => "000100110110010011", xin_1 => "000101001110111110", pass => true),
  (xin_0 => "000101111100001011", xin_1 => "001001110110100010", pass => false),
  (xin_0 => "000111011111011010", xin_1 => "001001110001011111", pass => false),
  (xin_0 => "001000010110101101", xin_1 => "000010000100001000", pass => false),
  (xin_0 => "001000010111001011", xin_1 => "000001100010010111", pass => false),
  (xin_0 => "001000010101010011", xin_1 => "001011000001110101", pass => false),
  (xin_0 => "001010111100100101", xin_1 => "000011100011101011", pass => true),
  (xin_0 => "001010000010000011", xin_1 => "001011000101101010", pass => false),
  (xin_0 => "001001001110001100", xin_1 => "000011001001000110", pass => false),
  (xin_0 => "001011100101001111", xin_1 => "000110110011110010", pass => false),
  (xin_0 => "001001110101001010", xin_1 => "000010000111001010", pass => false),
  (xin_0 => "001000100101111010", xin_1 => "000001101101111001", pass => false),
  (xin_0 => "001010100100011110", xin_1 => "000010111111100010", pass => true),
  (xin_0 => "001010101001110010", xin_1 => "000101010010000100", pass => true),
  (xin_0 => "001010000010111110", xin_1 => "000110110101001001", pass => true),
  (xin_0 => "001011010010001111", xin_1 => "001001111010011000", pass => false),
  (xin_0 => "000111001110101000", xin_1 => "001010101010100010", pass => false),
  (xin_0 => "001011001011011001", xin_1 => "000011010010101000", pass => true),
  (xin_0 => "001010111100000001", xin_1 => "001100111001111100", pass => false),
  (xin_0 => "001000100011010101", xin_1 => "000110000100011000", pass => true),
  (xin_0 => "001100110010111001", xin_1 => "000111001111110000", pass => false),
  (xin_0 => "001000100101110001", xin_1 => "000111110011111011", pass => true),
  (xin_0 => "001001100001011001", xin_1 => "000001000010110011", pass => false),
  (xin_0 => "000110010000101101", xin_1 => "000010000000110001", pass => false),
  (xin_0 => "001010011111101100", xin_1 => "000110000110001100", pass => true),
  (xin_0 => "001000000100011010", xin_1 => "001001110011100111", pass => false),
  (xin_0 => "001000000100101110", xin_1 => "001010110001101100", pass => false),
  (xin_0 => "001010110111010010", xin_1 => "001001011110101110", pass => false),
  (xin_0 => "001011010001101100", xin_1 => "001000110100010110", pass => false),
  (xin_0 => "000111101100100101", xin_1 => "001100001111011111", pass => false),
  (xin_0 => "000111110000011101", xin_1 => "000110011001010101", pass => true),
  (xin_0 => "000101010101111011", xin_1 => "001000110101010010", pass => false),
  (xin_0 => "001000100100100110", xin_1 => "000010000011110111", pass => false),
  (xin_0 => "000111001010001000", xin_1 => "000011111100111110", pass => false),
  (xin_0 => "001001100111100010", xin_1 => "001000000101110110", pass => true),
  (xin_0 => "000110110001011100", xin_1 => "000010111101000110", pass => false),
  (xin_0 => "001011000110011110", xin_1 => "000010100100111010", pass => true),
  (xin_0 => "001001010000011001", xin_1 => "000110100010100100", pass => true),
  (xin_0 => "001100010011000100", xin_1 => "000100110110110100", pass => true),
  (xin_0 => "001010001101000000", xin_1 => "000001011111100101", pass => false),
  (xin_0 => "000100100000101010", xin_1 => "001001111000111111", pass => false),
  (xin_0 => "000111010000101110", xin_1 => "001001010010111110", pass => false),
  (xin_0 => "001011001000100111", xin_1 => "001000100110100010", pass => false),
  (xin_0 => "001100001011110111", xin_1 => "000000111111100110", pass => true),
  (xin_0 => "001100011101011001", xin_1 => "000110111010110100", pass => false),
  (xin_0 => "001011110011101010", xin_1 => "000110100100101101", pass => false),
  (xin_0 => "001000110111011000", xin_1 => "001100101001010111", pass => false),
  (xin_0 => "001011100001010010", xin_1 => "000101010101101100", pass => true),
  (xin_0 => "001101001010101110", xin_1 => "001010010001111000", pass => true),
  (xin_0 => "010000101111101100", xin_1 => "001001100111111101", pass => true),
  (xin_0 => "000110100010011011", xin_1 => "001010100000001111", pass => false),
  (xin_0 => "000011111001010000", xin_1 => "000010010111010001", pass => true),
  (xin_0 => "001000101110111010", xin_1 => "000010110011101111", pass => false),
  (xin_0 => "000101001001100000", xin_1 => "001001000000110110", pass => false),
  (xin_0 => "000100000110001101", xin_1 => "001001000011011101", pass => false),
  (xin_0 => "001011100010000101", xin_1 => "001000110110101100", pass => false),
  (xin_0 => "001010101110111000", xin_1 => "001000111111001101", pass => false),
  (xin_0 => "000110111000011010", xin_1 => "000011010010000011", pass => false),
  (xin_0 => "000111011001111110", xin_1 => "000010011111101001", pass => false),
  (xin_0 => "001011010000000110", xin_1 => "001000110001001111", pass => false),
  (xin_0 => "001100101111010011", xin_1 => "000001000000010100", pass => true),
  (xin_0 => "000111111011000001", xin_1 => "000110000100100101", pass => true),
  (xin_0 => "001100001000001011", xin_1 => "001000011110100001", pass => false),
  (xin_0 => "000110110000000000", xin_1 => "000011100110111011", pass => false),
  (xin_0 => "001101100111111011", xin_1 => "001010011110001010", pass => true),
  (xin_0 => "001101000011010100", xin_1 => "001011001100010011", pass => true),
  (xin_0 => "000110011101000111", xin_1 => "001001010011000110", pass => false),
  (xin_0 => "001001101001001100", xin_1 => "001011100000111110", pass => false),
  (xin_0 => "000110110010011010", xin_1 => "000100000010100100", pass => false),
  (xin_0 => "000110011110110110", xin_1 => "000111010100001110", pass => true),
  (xin_0 => "000111001001111001", xin_1 => "000111100001010001", pass => true),
  (xin_0 => "001101101101010110", xin_1 => "000111110010010101", pass => false),
  (xin_0 => "001000111011110110", xin_1 => "001010111101111110", pass => false),
  (xin_0 => "000101101110100011", xin_1 => "000111100100000000", pass => true),
  (xin_0 => "000111001000011111", xin_1 => "001000000011100011", pass => true),
  (xin_0 => "000100101101001011", xin_1 => "000110000111100110", pass => true),
  (xin_0 => "001001110101001100", xin_1 => "000010101000001010", pass => false),
  (xin_0 => "000111001110010000", xin_1 => "000001010111110101", pass => false),
  (xin_0 => "001010001100001110", xin_1 => "001100010001110110", pass => false),
  (xin_0 => "000101111111010100", xin_1 => "000111011110000011", pass => true),
  (xin_0 => "001000000001001100", xin_1 => "000101011011010001", pass => true),
  (xin_0 => "001000100101101101", xin_1 => "000001001001001110", pass => false),
  (xin_0 => "000110111101011100", xin_1 => "001000011000100010", pass => true),
  (xin_0 => "001001110110100010", xin_1 => "000111111101011011", pass => true),
  (xin_0 => "000110010011100010", xin_1 => "000011011011101100", pass => false),
  (xin_0 => "000011100101001011", xin_1 => "000100110011100111", pass => true),
  (xin_0 => "001001000000001001", xin_1 => "000010100000010100", pass => false),
  (xin_0 => "001010111001110000", xin_1 => "001001011110001101", pass => false),
  (xin_0 => "000110011110101001", xin_1 => "000101000100111010", pass => true),
  (xin_0 => "001000010110000100", xin_1 => "000110101111110011", pass => true),
  (xin_0 => "001011110011111010", xin_1 => "001000110010011111", pass => false),
  (xin_0 => "000100010110011000", xin_1 => "000100001010010111", pass => true),
  (xin_0 => "001011011111001010", xin_1 => "000011111001000001", pass => true),
  (xin_0 => "001011000011010010", xin_1 => "000100011110111000", pass => true),
  (xin_0 => "000110100110100110", xin_1 => "000010101101111110", pass => false),
  (xin_0 => "000011100100011101", xin_1 => "000001110001000100", pass => true),
  (xin_0 => "001101111111111101", xin_1 => "001001001010000011", pass => true),
  (xin_0 => "000111000000110110", xin_1 => "000100100011100100", pass => true),
  (xin_0 => "000100110101111011", xin_1 => "000101001000100110", pass => true),
  (xin_0 => "001001110110000100", xin_1 => "000010001010010010", pass => false),
  (xin_0 => "001100101101001011", xin_1 => "000010010110000011", pass => true),
  (xin_0 => "000110001001100101", xin_1 => "000111010010010100", pass => true),
  (xin_0 => "000111111110111001", xin_1 => "000001000110011001", pass => false),
  (xin_0 => "001010001101011011", xin_1 => "001100111001011010", pass => false),
  (xin_0 => "001100000101011100", xin_1 => "001001000010011100", pass => false),
  (xin_0 => "000111110011111010", xin_1 => "001011000110100010", pass => false),
  (xin_0 => "000111100110010110", xin_1 => "000001101000101100", pass => false),
  (xin_0 => "001011111011011001", xin_1 => "001011000111010000", pass => false),
  (xin_0 => "001101001000101111", xin_1 => "001010011011111110", pass => true),
  (xin_0 => "001101001000111111", xin_1 => "000010011101111100", pass => true),
  (xin_0 => "001001111110010010", xin_1 => "000111001111010001", pass => true),
  (xin_0 => "001001000000110011", xin_1 => "001001111110011101", pass => false),
  (xin_0 => "000101100111101001", xin_1 => "000110000100111000", pass => true),
  (xin_0 => "001000101000110110", xin_1 => "000010011011011101", pass => false),
  (xin_0 => "001001111110000100", xin_1 => "000011010010111011", pass => false),
  (xin_0 => "001000001101111110", xin_1 => "000011011001010101", pass => false),
  (xin_0 => "000101110101110101", xin_1 => "000101010011000010", pass => true),
  (xin_0 => "000111111010010011", xin_1 => "000010010101101011", pass => false),
  (xin_0 => "001001111101111101", xin_1 => "001001111011110001", pass => false),
  (xin_0 => "001001110010110101", xin_1 => "000100110001000100", pass => true),
  (xin_0 => "001000001111111001", xin_1 => "000010011100100010", pass => false),
  (xin_0 => "000111101100101101", xin_1 => "000010110011010100", pass => false),
  (xin_0 => "000011011010101011", xin_1 => "111111011011101010", pass => true),
  (xin_0 => "000101110111100110", xin_1 => "000010011100110111", pass => false),
  (xin_0 => "001110100010010010", xin_1 => "001010100000011111", pass => true),
  (xin_0 => "000110001111100000", xin_1 => "000001101010101101", pass => false),
  (xin_0 => "001011100011010101", xin_1 => "000111000111110100", pass => false),
  (xin_0 => "000011101000110000", xin_1 => "000011111101011101", pass => true),
  (xin_0 => "001000011010100100", xin_1 => "000101111100100100", pass => true),
  (xin_0 => "001101101101001101", xin_1 => "000110010111110101", pass => false),
  (xin_0 => "001000000011100001", xin_1 => "000010000010110101", pass => false),
  (xin_0 => "001000111111000001", xin_1 => "000101000101000000", pass => true),
  (xin_0 => "000100100001110111", xin_1 => "000110101000001111", pass => true),
  (xin_0 => "000111110100100111", xin_1 => "000101100101111110", pass => true),
  (xin_0 => "001010111110011011", xin_1 => "001001010100111100", pass => false),
  (xin_0 => "000100110101100100", xin_1 => "001000011100001100", pass => false),
  (xin_0 => "000111001011001101", xin_1 => "000010100001101000", pass => false),
  (xin_0 => "000110110110110001", xin_1 => "000110111000011111", pass => true),
  (xin_0 => "000110111111011100", xin_1 => "000001111100111001", pass => false),
  (xin_0 => "001100001010001001", xin_1 => "000110110110011110", pass => false),
  (xin_0 => "000111010101011101", xin_1 => "000111111101111011", pass => true),
  (xin_0 => "001001001000111100", xin_1 => "000010010101000110", pass => false),
  (xin_0 => "000101101010111010", xin_1 => "000011000000010010", pass => false),
  (xin_0 => "001000001110101011", xin_1 => "000010011111001111", pass => false),
  (xin_0 => "001010011110111000", xin_1 => "000011000011110011", pass => true),
  (xin_0 => "000111101100010011", xin_1 => "000010111101001100", pass => false),
  (xin_0 => "000111101100111000", xin_1 => "000010001001011101", pass => false),
  (xin_0 => "001100110011110111", xin_1 => "000111011101100000", pass => false),
  (xin_0 => "000110101000110001", xin_1 => "001001100110110101", pass => false),
  (xin_0 => "000111101110111101", xin_1 => "000100000000011011", pass => false),
  (xin_0 => "000111111011011101", xin_1 => "000011101011111111", pass => false),
  (xin_0 => "001011110010001000", xin_1 => "001000000010110001", pass => false),
  (xin_0 => "001001101100110110", xin_1 => "000111001010101001", pass => true),
  (xin_0 => "000011010110110000", xin_1 => "000111110100110000", pass => false),
  (xin_0 => "001010110010000000", xin_1 => "000100001011011111", pass => true),
  (xin_0 => "000100101000001100", xin_1 => "000111111010100001", pass => false),
  (xin_0 => "001000110000101001", xin_1 => "000110011011010101", pass => true),
  (xin_0 => "001011111011001010", xin_1 => "000101000100001111", pass => true),
  (xin_0 => "000110110111011110", xin_1 => "000010000000001111", pass => false),
  (xin_0 => "001000101001101001", xin_1 => "000111101011111110", pass => true),
  (xin_0 => "001100000000000110", xin_1 => "001000001101010000", pass => false),
  (xin_0 => "001001110101001100", xin_1 => "000101110010110011", pass => true),
  (xin_0 => "000101111111101001", xin_1 => "000010101000000001", pass => false),
  (xin_0 => "001001010011100100", xin_1 => "001000000011001001", pass => true),
  (xin_0 => "000110101011110001", xin_1 => "001001000011101111", pass => false),
  (xin_0 => "001011000000010111", xin_1 => "001001001001100010", pass => false),
  (xin_0 => "000111000100000110", xin_1 => "000001100010001111", pass => false),
  (xin_0 => "001100010110011100", xin_1 => "000001111101111001", pass => true),
  (xin_0 => "000111011100001110", xin_1 => "000110110110101001", pass => true),
  (xin_0 => "001010010110010100", xin_1 => "000100001111011110", pass => true),
  (xin_0 => "001101100000101111", xin_1 => "001001110000001101", pass => true),
  (xin_0 => "001000101111110000", xin_1 => "001010100001010100", pass => false),
  (xin_0 => "000101100010101100", xin_1 => "000111100000101001", pass => true),
  (xin_0 => "001110011001011100", xin_1 => "000101110011001001", pass => false),
  (xin_0 => "001000110110100101", xin_1 => "001010001100000010", pass => false),
  (xin_0 => "001100011011101001", xin_1 => "000011010110000111", pass => true),
  (xin_0 => "000100111010011001", xin_1 => "000100110010011010", pass => true),
  (xin_0 => "001001000111010001", xin_1 => "000101110011011011", pass => true),
  (xin_0 => "001001000010010001", xin_1 => "001011001001100101", pass => false),
  (xin_0 => "000100011110111000", xin_1 => "000100010110011001", pass => true),
  (xin_0 => "001010110111110011", xin_1 => "001010101111111110", pass => false),
  (xin_0 => "001100110011111100", xin_1 => "000001000001100110", pass => true),
  (xin_0 => "001010010001101101", xin_1 => "000110110011110010", pass => true),
  (xin_0 => "001101010000011110", xin_1 => "000111010101100110", pass => false),
  (xin_0 => "000111100111000111", xin_1 => "000011001011000001", pass => false),
  (xin_0 => "000111011100011111", xin_1 => "001001111000100010", pass => false),
  (xin_0 => "001011110000111111", xin_1 => "001000001011000111", pass => false),
  (xin_0 => "001000100001100101", xin_1 => "000010000011110110", pass => false),
  (xin_0 => "000011100111010000", xin_1 => "000001001111001111", pass => true),
  (xin_0 => "000100011010001001", xin_1 => "000100100001100000", pass => true),
  (xin_0 => "000110010101111101", xin_1 => "000010110010110011", pass => false),
  (xin_0 => "000110001111100001", xin_1 => "001001010100011010", pass => false),
  (xin_0 => "000111000111011000", xin_1 => "001001100001001000", pass => false),
  (xin_0 => "001000111000100110", xin_1 => "000111001001011111", pass => true),
  (xin_0 => "001101000010001111", xin_1 => "000011110001011000", pass => true),
  (xin_0 => "000110011101010111", xin_1 => "000010100011100101", pass => false),
  (xin_0 => "000110100011111100", xin_1 => "000111101100001001", pass => true),
  (xin_0 => "001011111010100000", xin_1 => "001001001100011001", pass => false),
  (xin_0 => "001100110111011010", xin_1 => "000001101001010011", pass => true),
  (xin_0 => "000101110010001001", xin_1 => "000111000110110000", pass => true),
  (xin_0 => "001000010101010101", xin_1 => "000111011000011100", pass => true),
  (xin_0 => "000110010001101011", xin_1 => "000101111010101011", pass => true),
  (xin_0 => "000110011100100101", xin_1 => "001011000100111101", pass => false),
  (xin_0 => "000111000010000000", xin_1 => "000001110000101010", pass => false),
  (xin_0 => "000100001110001001", xin_1 => "000101001000000010", pass => true),
  (xin_0 => "000101101001111000", xin_1 => "001001100001000000", pass => false),
  (xin_0 => "000011000001110100", xin_1 => "000110101000000000", pass => false),
  (xin_0 => "000110101111011010", xin_1 => "000110111000111001", pass => true),
  (xin_0 => "001100001111100101", xin_1 => "000101111000011011", pass => false),
  (xin_0 => "001000000110010000", xin_1 => "000010010111001001", pass => false),
  (xin_0 => "001110000011111101", xin_1 => "001010101110111100", pass => true),
  (xin_0 => "000101110001110000", xin_1 => "000110101000110101", pass => true),
  (xin_0 => "001011101000100101", xin_1 => "001000111100101111", pass => false),
  (xin_0 => "000111110000101110", xin_1 => "000010001001011011", pass => false),
  (xin_0 => "001001000011110101", xin_1 => "000101100000000010", pass => true),
  (xin_0 => "001001001110111001", xin_1 => "000010111000001011", pass => false),
  (xin_0 => "001100101101010000", xin_1 => "000110001001000111", pass => false),
  (xin_0 => "001010010001100111", xin_1 => "000111000100100110", pass => true),
  (xin_0 => "000101111000001101", xin_1 => "001001000001000001", pass => false),
  (xin_0 => "000110111101101000", xin_1 => "000010010100100011", pass => false),
  (xin_0 => "001000000101100100", xin_1 => "000001111101110110", pass => false),
  (xin_0 => "000100110100110101", xin_1 => "000001101000001111", pass => true),
  (xin_0 => "001100010000011011", xin_1 => "000011010111111111", pass => true),
  (xin_0 => "000110111001100010", xin_1 => "000101011011100110", pass => true),
  (xin_0 => "000110101010001010", xin_1 => "000101110100110111", pass => true),
  (xin_0 => "001101110001000110", xin_1 => "001010100010011001", pass => true),
  (xin_0 => "001000110111011101", xin_1 => "001000000110100011", pass => true),
  (xin_0 => "001010001100010100", xin_1 => "000001111000011111", pass => false),
  (xin_0 => "001010110000101100", xin_1 => "001001100100110100", pass => false),
  (xin_0 => "000101011110100011", xin_1 => "000100110110111001", pass => true),
  (xin_0 => "001011110100100011", xin_1 => "000101111111101111", pass => true),
  (xin_0 => "001110100111101000", xin_1 => "001010000111111100", pass => true),
  (xin_0 => "001010101110010000", xin_1 => "001001001100110110", pass => false),
  (xin_0 => "000110000110101111", xin_1 => "001001011101001110", pass => false),
  (xin_0 => "001100001101001000", xin_1 => "001000001000010001", pass => false),
  (xin_0 => "001001010101000100", xin_1 => "001010100001011010", pass => false),
  (xin_0 => "001100101111001001", xin_1 => "000101001000011111", pass => true),
  (xin_0 => "000111011000000010", xin_1 => "000011111000000110", pass => false),
  (xin_0 => "000110010111011100", xin_1 => "000010011000011100", pass => false),
  (xin_0 => "001001000100000101", xin_1 => "000110101111000011", pass => true),
  (xin_0 => "001010001111100110", xin_1 => "000110010111111111", pass => true),
  (xin_0 => "000111111100100101", xin_1 => "000100100010011000", pass => true),
  (xin_0 => "001011101101011110", xin_1 => "001000110001010010", pass => false),
  (xin_0 => "001001000010110001", xin_1 => "000011010000010101", pass => false),
  (xin_0 => "001100011101110000", xin_1 => "000011110111111101", pass => true),
  (xin_0 => "000111110001001001", xin_1 => "000111010010011001", pass => true),
  (xin_0 => "000011001011000111", xin_1 => "000111111001011001", pass => false),
  (xin_0 => "001011001011001010", xin_1 => "000101011110011010", pass => true),
  (xin_0 => "000110011100011010", xin_1 => "000101101000010011", pass => true),
  (xin_0 => "001000010000111000", xin_1 => "000110100111000011", pass => true),
  (xin_0 => "001000010100010000", xin_1 => "000010000001110111", pass => false),
  (xin_0 => "001011101000101011", xin_1 => "000010101010101001", pass => true),
  (xin_0 => "001100100010101011", xin_1 => "001000101000001100", pass => false),
  (xin_0 => "001100000110001001", xin_1 => "000011001100101110", pass => true),
  (xin_0 => "000101111001111101", xin_1 => "000011101100101000", pass => true),
  (xin_0 => "001011111010000010", xin_1 => "000101011011101111", pass => true),
  (xin_0 => "000111011000000111", xin_1 => "000011101100111111", pass => false),
  (xin_0 => "000110001001110111", xin_1 => "000100010100011110", pass => true),
  (xin_0 => "001100010010010100", xin_1 => "001000011001101101", pass => false),
  (xin_0 => "001001001001000110", xin_1 => "000011111001100111", pass => false),
  (xin_0 => "001000010101111001", xin_1 => "000100101110111011", pass => true),
  (xin_0 => "000101001111111100", xin_1 => "000110110111111011", pass => true),
  (xin_0 => "001011010001001111", xin_1 => "001001010000000100", pass => false),
  (xin_0 => "001010100000001000", xin_1 => "001100010001111010", pass => false),
  (xin_0 => "000110100100011000", xin_1 => "001000011100011101", pass => false),
  (xin_0 => "000110101101111001", xin_1 => "001001000100000100", pass => false),
  (xin_0 => "001001110011011100", xin_1 => "000001101011010010", pass => false),
  (xin_0 => "000110111111101101", xin_1 => "001010001011100100", pass => false),
  (xin_0 => "001010011111001011", xin_1 => "001011001001001011", pass => false),
  (xin_0 => "000111011111000101", xin_1 => "000111010011111101", pass => true),
  (xin_0 => "000011010010111011", xin_1 => "000011011111100001", pass => true),
  (xin_0 => "000111010111000100", xin_1 => "000010111110001100", pass => false),
  (xin_0 => "000110100011110111", xin_1 => "000001001000111001", pass => false),
  (xin_0 => "001001100101101111", xin_1 => "001100100011011001", pass => false),
  (xin_0 => "000100010101011101", xin_1 => "000010000110100110", pass => true),
  (xin_0 => "000110001010000100", xin_1 => "000011010000001111", pass => false),
  (xin_0 => "001100011111011100", xin_1 => "001010101110001010", pass => true),
  (xin_0 => "000111110110101100", xin_1 => "001000001010101110", pass => true),
  (xin_0 => "001000000010100011", xin_1 => "000010111001101011", pass => false),
  (xin_0 => "001000011111100110", xin_1 => "000101110111010000", pass => true),
  (xin_0 => "000101011110010100", xin_1 => "000101011110001110", pass => true),
  (xin_0 => "001011000001000011", xin_1 => "001000110001011011", pass => false),
  (xin_0 => "000111010010110001", xin_1 => "000011100011011011", pass => false),
  (xin_0 => "000100011100001001", xin_1 => "000101001110101001", pass => true),
  (xin_0 => "000011010111001111", xin_1 => "000101111101111001", pass => true),
  (xin_0 => "001100000111010100", xin_1 => "001001111010011111", pass => false),
  (xin_0 => "001011101000110001", xin_1 => "001001001011101101", pass => false),
  (xin_0 => "000111101001100000", xin_1 => "000001011001010111", pass => false),
  (xin_0 => "001101001011011000", xin_1 => "000011011101011111", pass => true),
  (xin_0 => "000110100101100001", xin_1 => "000010110110110100", pass => false),
  (xin_0 => "001011000111001011", xin_1 => "001000111001001100", pass => false),
  (xin_0 => "001011111010000000", xin_1 => "001000011100011011", pass => false),
  (xin_0 => "000101110101010000", xin_1 => "000100010111011101", pass => true),
  (xin_0 => "001101100100001110", xin_1 => "000100101000111101", pass => false),
  (xin_0 => "001001111001011010", xin_1 => "001010101000010111", pass => false),
  (xin_0 => "001011111000000010", xin_1 => "000111101011111010", pass => false),
  (xin_0 => "001001011010011010", xin_1 => "001010110011111110", pass => false),
  (xin_0 => "000111010100001110", xin_1 => "000011101000101011", pass => false),
  (xin_0 => "000011101011010100", xin_1 => "000111101010110001", pass => false),
  (xin_0 => "000110001101111000", xin_1 => "001001010100100010", pass => false),
  (xin_0 => "001110111101010101", xin_1 => "001001010101111000", pass => true),
  (xin_0 => "001000111101100001", xin_1 => "000110000011110001", pass => true),
  (xin_0 => "000111011111001010", xin_1 => "000010100100010001", pass => false),
  (xin_0 => "000101101110101000", xin_1 => "000100001111100010", pass => true),
  (xin_0 => "001100111011101001", xin_1 => "001001111111000011", pass => true),
  (xin_0 => "001011111111101100", xin_1 => "000111100110100111", pass => false),
  (xin_0 => "001100000000001111", xin_1 => "000111101010010011", pass => false),
  (xin_0 => "001010100110100011", xin_1 => "001001101101110100", pass => false),
  (xin_0 => "001000011110001011", xin_1 => "000110101110101110", pass => true),
  (xin_0 => "001000110000000000", xin_1 => "000010011111111001", pass => false),
  (xin_0 => "001100001111011110", xin_1 => "000111100001111110", pass => false),
  (xin_0 => "000100101110100001", xin_1 => "000011100001010100", pass => true),
  (xin_0 => "001100011000001011", xin_1 => "000110011110001000", pass => false),
  (xin_0 => "000110100001101011", xin_1 => "001000001011110111", pass => true),
  (xin_0 => "001101101011111011", xin_1 => "000110011001001010", pass => false),
  (xin_0 => "000111111101000001", xin_1 => "000111010111110000", pass => true),
  (xin_0 => "000010111000000111", xin_1 => "000011000001000110", pass => true),
  (xin_0 => "001010101101000011", xin_1 => "000111111010100011", pass => false),
  (xin_0 => "000011101010110011", xin_1 => "000100001101001100", pass => true),
  (xin_0 => "001010001101001010", xin_1 => "001000100000010100", pass => false),
  (xin_0 => "001001011000111011", xin_1 => "000111001101000111", pass => true),
  (xin_0 => "001101001011011100", xin_1 => "000100101011100110", pass => true),
  (xin_0 => "001101011011000101", xin_1 => "001010000000100111", pass => true),
  (xin_0 => "000100010111100111", xin_1 => "001000101011100101", pass => false),
  (xin_0 => "000101110000110101", xin_1 => "001000101101100000", pass => false),
  (xin_0 => "001010001000000110", xin_1 => "000010100101000010", pass => false),
  (xin_0 => "000101100001011101", xin_1 => "000011011111110111", pass => true),
  (xin_0 => "001011000101000001", xin_1 => "001001000010110000", pass => false),
  (xin_0 => "000011100011011100", xin_1 => "000000110100011110", pass => true),
  (xin_0 => "001000010011100101", xin_1 => "000100111100111110", pass => true),
  (xin_0 => "001110101010010100", xin_1 => "001001001111001110", pass => true),
  (xin_0 => "001001100001011001", xin_1 => "000011110111000111", pass => false),
  (xin_0 => "001000110110001101", xin_1 => "000101110010100010", pass => true),
  (xin_0 => "000110111000010100", xin_1 => "000001101101010000", pass => false),
  (xin_0 => "000101111011111111", xin_1 => "000010111101000110", pass => false),
  (xin_0 => "001100111010011101", xin_1 => "000110111001001011", pass => false),
  (xin_0 => "000110111111001000", xin_1 => "000101111011111100", pass => true),
  (xin_0 => "001001111010010010", xin_1 => "000001101110000110", pass => false),
  (xin_0 => "001000101001011011", xin_1 => "000101010001001000", pass => true),
  (xin_0 => "001011001010011100", xin_1 => "001001000001101101", pass => false),
  (xin_0 => "001100011101110100", xin_1 => "000110101011111101", pass => false),
  (xin_0 => "000110111001111100", xin_1 => "000001111000011101", pass => false),
  (xin_0 => "000111000001011001", xin_1 => "000011100000011000", pass => false),
  (xin_0 => "001001001111110000", xin_1 => "000010000000101110", pass => false),
  (xin_0 => "001010100011010101", xin_1 => "001001001001100100", pass => false),
  (xin_0 => "000101001000011011", xin_1 => "001001100100001100", pass => false),
  (xin_0 => "000001011010110010", xin_1 => "000110111000101111", pass => false),
  (xin_0 => "000110001101001010", xin_1 => "000011001111011100", pass => false),
  (xin_0 => "001001110000001100", xin_1 => "000111011011111000", pass => true),
  (xin_0 => "001001010000011001", xin_1 => "000001001001100011", pass => false),
  (xin_0 => "001011111100000010", xin_1 => "000010110100000111", pass => true),
  (xin_0 => "001111001110110101", xin_1 => "001010101000010101", pass => true),
  (xin_0 => "001100000100101001", xin_1 => "000000101010000011", pass => true),
  (xin_0 => "001000110100110111", xin_1 => "000111001001111101", pass => true),
  (xin_0 => "000111000000011100", xin_1 => "001010010101001111", pass => false),
  (xin_0 => "001011011001100011", xin_1 => "000110111101110001", pass => false),
  (xin_0 => "001010111011100101", xin_1 => "001001011110000001", pass => false),
  (xin_0 => "000101110110111000", xin_1 => "000110001111100100", pass => true),
  (xin_0 => "001100010100001100", xin_1 => "001001001100110101", pass => false),
  (xin_0 => "000110110001100111", xin_1 => "000101110111110100", pass => true),
  (xin_0 => "000011010100100100", xin_1 => "001000110000011011", pass => false),
  (xin_0 => "000101101011110111", xin_1 => "000100111000011010", pass => true),
  (xin_0 => "001100011010100011", xin_1 => "000110100100111000", pass => false),
  (xin_0 => "000101100001001000", xin_1 => "001001010011000111", pass => false),
  (xin_0 => "000011110100101101", xin_1 => "000010100111010111", pass => true),
  (xin_0 => "000011001011110011", xin_1 => "000011011101001000", pass => true),
  (xin_0 => "001011011101101011", xin_1 => "000011011100000100", pass => true),
  (xin_0 => "000100001110001110", xin_1 => "000001111011010101", pass => true),
  (xin_0 => "000011000000011011", xin_1 => "000001111101111100", pass => true),
  (xin_0 => "001110001111100100", xin_1 => "000111010010011001", pass => false),
  (xin_0 => "001001101010000000", xin_1 => "000111001001110001", pass => true),
  (xin_0 => "001001101001000001", xin_1 => "000110010101101101", pass => true),
  (xin_0 => "000100010011111010", xin_1 => "001000100111111001", pass => false),
  (xin_0 => "000111111011101110", xin_1 => "000100101111001111", pass => true),
  (xin_0 => "001110100111100111", xin_1 => "001010001100111101", pass => true),
  (xin_0 => "001100100011011110", xin_1 => "000010001011011110", pass => true),
  (xin_0 => "001000110000011100", xin_1 => "001011100000010010", pass => false),
  (xin_0 => "001011100101010011", xin_1 => "000110100111010101", pass => false),
  (xin_0 => "001000110001101011", xin_1 => "000001111110000011", pass => false),
  (xin_0 => "001110011110100001", xin_1 => "001010011001001010", pass => true),
  (xin_0 => "001001011011101010", xin_1 => "000001011011010111", pass => false),
  (xin_0 => "001010010000100010", xin_1 => "001011000110001011", pass => false),
  (xin_0 => "000100001111111011", xin_1 => "000110110111111110", pass => false),
  (xin_0 => "000100111110010100", xin_1 => "000101110110100011", pass => true),
  (xin_0 => "001011000001110000", xin_1 => "000111101101010101", pass => false),
  (xin_0 => "001101110101010111", xin_1 => "000100110010101010", pass => false),
  (xin_0 => "000100011001000111", xin_1 => "001000010010100111", pass => false),
  (xin_0 => "001000110011000011", xin_1 => "000001100111011110", pass => false),
  (xin_0 => "000111000100010101", xin_1 => "000101101111101100", pass => true),
  (xin_0 => "001001011001111000", xin_1 => "000110101100001101", pass => true),
  (xin_0 => "001011011010010110", xin_1 => "000111011100110000", pass => false),
  (xin_0 => "001100001101001010", xin_1 => "001000110110001101", pass => false),
  (xin_0 => "000111001111111100", xin_1 => "000010001000101101", pass => false),
  (xin_0 => "001100000111101011", xin_1 => "000010011110000001", pass => true),
  (xin_0 => "000110001000011110", xin_1 => "000111101110111011", pass => true),
  (xin_0 => "001011010011100100", xin_1 => "000101101000100101", pass => true),
  (xin_0 => "001100100000101000", xin_1 => "000101111011001010", pass => false),
  (xin_0 => "000111001011111001", xin_1 => "000110010000010010", pass => true),
  (xin_0 => "001100110011111110", xin_1 => "000101111110111101", pass => false),
  (xin_0 => "001010111010011100", xin_1 => "001000111100000001", pass => false),
  (xin_0 => "001010011011010000", xin_1 => "000101001110001000", pass => true),
  (xin_0 => "001010110100001010", xin_1 => "000101000000000111", pass => true),
  (xin_0 => "000100111001010011", xin_1 => "000111000001010001", pass => true),
  (xin_0 => "001011010111001111", xin_1 => "001010010000110110", pass => false),
  (xin_0 => "000011101101110000", xin_1 => "000100010001100010", pass => true),
  (xin_0 => "000110001111001011", xin_1 => "000101111101110101", pass => true),
  (xin_0 => "000111000110100010", xin_1 => "000010000011001000", pass => false),
  (xin_0 => "001001010110110011", xin_1 => "000011001010100110", pass => false),
  (xin_0 => "000110011101010101", xin_1 => "000011010001011111", pass => false),
  (xin_0 => "001000010111100101", xin_1 => "001000011001000011", pass => true),
  (xin_0 => "001101001010001101", xin_1 => "000111000011101001", pass => false),
  (xin_0 => "001011010011010101", xin_1 => "000110010000010101", pass => true),
  (xin_0 => "001001000000100000", xin_1 => "000110011000100001", pass => true),
  (xin_0 => "010000001001100110", xin_1 => "001001111001001011", pass => true),
  (xin_0 => "001011000010111000", xin_1 => "000011010000110010", pass => true),
  (xin_0 => "000101110111101101", xin_1 => "000011100111010101", pass => true),
  (xin_0 => "000100000110101001", xin_1 => "001000111001101100", pass => false),
  (xin_0 => "000110001011001011", xin_1 => "001001100000000000", pass => false),
  (xin_0 => "001100010101100001", xin_1 => "001010011000011000", pass => false),
  (xin_0 => "001011110011010010", xin_1 => "000010001111011101", pass => true),
  (xin_0 => "001001011010101001", xin_1 => "000110110011010000", pass => true),
  (xin_0 => "001001000000001010", xin_1 => "000010011001110010", pass => false),
  (xin_0 => "001011011001110000", xin_1 => "001000100011101011", pass => false),
  (xin_0 => "001101000100010110", xin_1 => "001011101101011010", pass => true),
  (xin_0 => "001010100011011101", xin_1 => "001001011001011110", pass => false),
  (xin_0 => "001100000111110111", xin_1 => "001001010110001110", pass => false),
  (xin_0 => "000101000100001000", xin_1 => "000100110100100110", pass => true),
  (xin_0 => "000110101110100011", xin_1 => "000011011101101011", pass => false),
  (xin_0 => "000110110101110011", xin_1 => "001010011000101111", pass => false),
  (xin_0 => "000110101101000111", xin_1 => "000010011001111110", pass => false),
  (xin_0 => "000110110101111010", xin_1 => "001010110001011100", pass => false),
  (xin_0 => "001001001010100011", xin_1 => "000110001110001111", pass => true),
  (xin_0 => "000111110110100110", xin_1 => "000010011000010111", pass => false),
  (xin_0 => "010000101101110101", xin_1 => "001001110010011000", pass => true),
  (xin_0 => "001000001100000110", xin_1 => "000010110001011100", pass => false),
  (xin_0 => "000111101100011100", xin_1 => "000010101100001010", pass => false),
  (xin_0 => "001001000011011010", xin_1 => "000100001000001100", pass => false),
  (xin_0 => "000110110001100001", xin_1 => "000111010001000001", pass => true),
  (xin_0 => "001010100001101100", xin_1 => "001001000000001100", pass => false),
  (xin_0 => "001110011000110010", xin_1 => "000101010110010000", pass => false),
  (xin_0 => "000111110000100111", xin_1 => "000111101110010111", pass => true),
  (xin_0 => "001001010101000011", xin_1 => "000100110011010110", pass => true),
  (xin_0 => "000111000111000011", xin_1 => "001010010100101101", pass => false),
  (xin_0 => "000011100001111010", xin_1 => "000010001101101001", pass => true),
  (xin_0 => "001101010011011101", xin_1 => "000111110111101110", pass => false),
  (xin_0 => "010000001110010011", xin_1 => "001001100110001111", pass => true),
  (xin_0 => "001100010111111001", xin_1 => "000110000100100101", pass => false),
  (xin_0 => "000101000100101001", xin_1 => "001000110111100010", pass => false),
  (xin_0 => "001001111000011000", xin_1 => "000100110100001100", pass => true),
  (xin_0 => "001110101010101000", xin_1 => "000110010110100010", pass => false),
  (xin_0 => "000111100101011100", xin_1 => "000010101101011000", pass => false),
  (xin_0 => "001100001101100010", xin_1 => "000011011101111000", pass => true),
  (xin_0 => "001010001010010100", xin_1 => "000111010010010110", pass => true),
  (xin_0 => "000110010100110011", xin_1 => "000111011111100001", pass => true),
  (xin_0 => "000101111111011000", xin_1 => "001001001010110100", pass => false),
  (xin_0 => "000110011001100101", xin_1 => "000001011001001011", pass => false),
  (xin_0 => "000110110111111110", xin_1 => "001001010010000010", pass => false),
  (xin_0 => "001011100010101101", xin_1 => "000101001110111101", pass => true),
  (xin_0 => "001001111100101101", xin_1 => "000010110001001110", pass => false),
  (xin_0 => "001100101001001100", xin_1 => "000100001011001110", pass => true),
  (xin_0 => "000100000011100110", xin_1 => "001000010111111100", pass => false),
  (xin_0 => "000111101001011011", xin_1 => "001000100101011000", pass => true),
  (xin_0 => "001100011011001101", xin_1 => "000110011100000001", pass => false),
  (xin_0 => "001000110110110000", xin_1 => "000010000101001001", pass => false),
  (xin_0 => "000100111110000111", xin_1 => "000101100110101100", pass => true),
  (xin_0 => "000110010110101001", xin_1 => "000011010001100010", pass => false),
  (xin_0 => "001101101001101101", xin_1 => "001001110110000000", pass => true),
  (xin_0 => "001000011100111101", xin_1 => "001011000100101110", pass => false),
  (xin_0 => "000110100111111110", xin_1 => "000111011011101010", pass => true),
  (xin_0 => "001000010001110100", xin_1 => "001000000001111100", pass => true),
  (xin_0 => "000110101110100110", xin_1 => "000110001011010101", pass => true),
  (xin_0 => "001000010110000010", xin_1 => "001010010100110010", pass => false),
  (xin_0 => "000100110110111111", xin_1 => "001001101101010011", pass => false),
  (xin_0 => "001000101101001100", xin_1 => "000010110100100000", pass => false),
  (xin_0 => "000110000000100010", xin_1 => "000101010101000100", pass => true),
  (xin_0 => "001000101011010001", xin_1 => "000011000001010100", pass => false),
  (xin_0 => "001001101000110000", xin_1 => "000111100100101100", pass => true),
  (xin_0 => "001101000011101110", xin_1 => "000110000101100001", pass => false),
  (xin_0 => "000100010010001110", xin_1 => "000010110010011101", pass => true),
  (xin_0 => "000110001000010001", xin_1 => "000101101011000100", pass => true),
  (xin_0 => "000111101100000101", xin_1 => "001000101110001101", pass => true),
  (xin_0 => "000101000110010010", xin_1 => "000101000010010011", pass => true),
  (xin_0 => "000111010001011001", xin_1 => "001010010011110101", pass => false),
  (xin_0 => "001001000110000101", xin_1 => "000010000101001001", pass => false),
  (xin_0 => "000010111000100000", xin_1 => "001000000100000010", pass => false),
  (xin_0 => "001101000101101000", xin_1 => "000011101111110000", pass => true),
  (xin_0 => "001100101111000001", xin_1 => "000001111110000101", pass => true),
  (xin_0 => "000011001001100111", xin_1 => "111111110110101110", pass => true),
  (xin_0 => "000110011110100010", xin_1 => "001001111011110111", pass => false),
  (xin_0 => "000110000010001000", xin_1 => "000001100100010001", pass => false),
  (xin_0 => "001100001101000101", xin_1 => "001000101110011001", pass => false),
  (xin_0 => "001010000011000110", xin_1 => "000100100001101001", pass => true),
  (xin_0 => "001011100011101011", xin_1 => "000101100000111001", pass => true),
  (xin_0 => "000110111101100100", xin_1 => "001001010011011101", pass => false),
  (xin_0 => "000110101011101010", xin_1 => "001001001011000000", pass => false),
  (xin_0 => "000100100010100011", xin_1 => "000111011010000000", pass => false),
  (xin_0 => "000110100000100010", xin_1 => "000111010110101100", pass => true),
  (xin_0 => "001101111010010111", xin_1 => "000100111100000011", pass => false),
  (xin_0 => "001001110001010010", xin_1 => "000011111010100001", pass => true),
  (xin_0 => "001011100010101010", xin_1 => "000111010001101000", pass => false),
  (xin_0 => "001000100001010111", xin_1 => "001000101101001110", pass => true),
  (xin_0 => "001010001001111111", xin_1 => "001001001110011110", pass => false),
  (xin_0 => "000111111010101110", xin_1 => "001010110011110100", pass => false),
  (xin_0 => "001010000001010010", xin_1 => "000011101000000101", pass => false),
  (xin_0 => "000101100010100100", xin_1 => "001001110010001001", pass => false),
  (xin_0 => "001110010100111001", xin_1 => "001010011010010010", pass => true),
  (xin_0 => "000100101111000011", xin_1 => "000101101011110100", pass => true),
  (xin_0 => "001110011110001001", xin_1 => "001010000101011000", pass => true),
  (xin_0 => "001100101101110111", xin_1 => "000111111010100011", pass => false),
  (xin_0 => "001010110000101100", xin_1 => "001000000111011010", pass => false),
  (xin_0 => "000111010011110010", xin_1 => "000010101111111100", pass => false),
  (xin_0 => "001111110000010100", xin_1 => "001001101011101000", pass => true),
  (xin_0 => "000101010101101000", xin_1 => "001001001110001000", pass => false),
  (xin_0 => "000011100100110001", xin_1 => "000001011101000110", pass => true),
  (xin_0 => "000101111101010000", xin_1 => "001001010010011011", pass => false),
  (xin_0 => "001011111000000010", xin_1 => "000011001111001001", pass => true),
  (xin_0 => "001011111101111011", xin_1 => "000111111100000010", pass => false),
  (xin_0 => "001000001111001111", xin_1 => "001000100101010011", pass => true),
  (xin_0 => "001100011111101011", xin_1 => "000110000101011111", pass => false),
  (xin_0 => "001011111101111011", xin_1 => "000010101010000111", pass => true),
  (xin_0 => "000110111000010000", xin_1 => "000010100110110111", pass => false),
  (xin_0 => "001000001100110000", xin_1 => "000010011110100011", pass => false),
  (xin_0 => "001101010111001101", xin_1 => "000010110011111001", pass => true),
  (xin_0 => "000110000100111101", xin_1 => "000110001011100010", pass => true),
  (xin_0 => "001001101001000111", xin_1 => "000001101000101111", pass => false),
  (xin_0 => "001100000101111111", xin_1 => "000110011111101100", pass => false),
  (xin_0 => "001100110000100111", xin_1 => "001001011110011101", pass => false),
  (xin_0 => "000110000101001011", xin_1 => "000110100100110000", pass => true),
  (xin_0 => "001000101011001111", xin_1 => "000001001011001100", pass => false),
  (xin_0 => "001001100111011011", xin_1 => "001011001011010011", pass => false),
  (xin_0 => "001000000100000010", xin_1 => "001001000101000110", pass => false),
  (xin_0 => "000111010001010101", xin_1 => "000101101011000101", pass => true),
  (xin_0 => "001001100101110110", xin_1 => "000011100101111101", pass => false),
  (xin_0 => "000101010101111100", xin_1 => "000100001110110111", pass => true),
  (xin_0 => "001100001010101010", xin_1 => "000111100010100000", pass => false),
  (xin_0 => "001011000010100011", xin_1 => "001000010010010111", pass => false),
  (xin_0 => "000111101011010100", xin_1 => "000001110100001111", pass => false),
  (xin_0 => "000110010110000000", xin_1 => "000001000111001000", pass => false),
  (xin_0 => "001001011111000110", xin_1 => "000111111011001011", pass => true),
  (xin_0 => "001000100011111010", xin_1 => "000010111000011011", pass => false),
  (xin_0 => "001001010001110000", xin_1 => "000110010100000111", pass => true),
  (xin_0 => "001001110110011001", xin_1 => "000100001000100101", pass => true),
  (xin_0 => "000110110001010100", xin_1 => "000010011011010001", pass => false),
  (xin_0 => "001100010101110110", xin_1 => "000111110001111001", pass => false),
  (xin_0 => "000111000001011010", xin_1 => "000010110111101111", pass => false),
  (xin_0 => "001000111001100101", xin_1 => "000010110010010111", pass => false),
  (xin_0 => "000110100111010100", xin_1 => "001001100111110010", pass => false),
  (xin_0 => "001000001111101000", xin_1 => "000010101001111000", pass => false),
  (xin_0 => "001100011000011101", xin_1 => "001000000010101110", pass => false),
  (xin_0 => "001011000011010000", xin_1 => "000111011111101011", pass => false),
  (xin_0 => "001000001101110011", xin_1 => "000101110010111100", pass => true),
  (xin_0 => "001100011001011111", xin_1 => "000111001010110001", pass => false),
  (xin_0 => "001010111010010000", xin_1 => "001000111010111100", pass => false),
  (xin_0 => "001101100111101001", xin_1 => "000111111111110001", pass => false),
  (xin_0 => "000111110101101111", xin_1 => "000010111100010111", pass => false),
  (xin_0 => "001011110101101111", xin_1 => "000110111010010001", pass => false),
  (xin_0 => "001100100011101001", xin_1 => "000101110010010001", pass => false),
  (xin_0 => "000110001011101000", xin_1 => "001001010001011101", pass => false),
  (xin_0 => "000110001000100000", xin_1 => "000101110110000011", pass => true),
  (xin_0 => "000111011100111010", xin_1 => "000011011100101100", pass => false),
  (xin_0 => "000110110011011010", xin_1 => "000111010100100101", pass => true),
  (xin_0 => "001001001110101001", xin_1 => "000010000000101101", pass => false),
  (xin_0 => "000111011001000101", xin_1 => "000010100011000110", pass => false),
  (xin_0 => "000101011010110010", xin_1 => "001001101000010100", pass => false),
  (xin_0 => "001000100010010000", xin_1 => "000011000110011001", pass => false),
  (xin_0 => "000100110000110011", xin_1 => "000110000001000000", pass => true),
  (xin_0 => "000110011101101000", xin_1 => "001010000010111011", pass => false),
  (xin_0 => "001010001110000111", xin_1 => "001101010111010100", pass => false),
  (xin_0 => "000011100100110001", xin_1 => "000011010011001100", pass => true),
  (xin_0 => "001011000011100001", xin_1 => "001010010000011011", pass => false),
  (xin_0 => "001010011100011110", xin_1 => "001000111010011111", pass => false),
  (xin_0 => "001100111001101001", xin_1 => "000100000000000101", pass => true),
  (xin_0 => "000111110000000001", xin_1 => "000010010010011100", pass => false),
  (xin_0 => "001000100100000001", xin_1 => "000110011100010100", pass => true),
  (xin_0 => "000111100110010101", xin_1 => "001010001011100001", pass => false),
  (xin_0 => "001000100100000100", xin_1 => "000010111001010010", pass => false),
  (xin_0 => "000100010110100111", xin_1 => "000011001011010010", pass => true),
  (xin_0 => "000110001101100111", xin_1 => "000101101000001111", pass => true),
  (xin_0 => "001011110010110011", xin_1 => "001000100011100011", pass => false),
  (xin_0 => "000101010110011000", xin_1 => "000110100010000001", pass => true),
  (xin_0 => "001001110101110010", xin_1 => "000010110001110001", pass => false),
  (xin_0 => "000111001011000010", xin_1 => "000010000101011001", pass => false),
  (xin_0 => "001101101101101000", xin_1 => "000101010010101001", pass => false),
  (xin_0 => "001001010111111100", xin_1 => "000100010100101110", pass => true),
  (xin_0 => "001100011101001100", xin_1 => "000111010011011011", pass => false),
  (xin_0 => "000110011100111011", xin_1 => "000111101111000111", pass => true),
  (xin_0 => "001010100101100001", xin_1 => "000010110010101001", pass => true),
  (xin_0 => "000011101001000101", xin_1 => "001000000011100011", pass => false),
  (xin_0 => "001010111100001100", xin_1 => "000101101001100111", pass => true),
  (xin_0 => "001011100111100111", xin_1 => "000100000011000011", pass => true),
  (xin_0 => "001010010111001101", xin_1 => "000110111110001011", pass => true),
  (xin_0 => "001010100010001100", xin_1 => "000010110100110100", pass => false),
  (xin_0 => "001001000010111010", xin_1 => "001010011100110101", pass => false),
  (xin_0 => "001010100001110101", xin_1 => "001001111100001010", pass => false),
  (xin_0 => "001100000010101011", xin_1 => "000111110010001110", pass => false),
  (xin_0 => "000110100101001110", xin_1 => "000011010111000110", pass => false),
  (xin_0 => "000101110100110000", xin_1 => "001001001110111010", pass => false),
  (xin_0 => "001001101100001011", xin_1 => "001101100110000110", pass => false),
  (xin_0 => "000110110010110111", xin_1 => "001001001110100101", pass => false),
  (xin_0 => "000100100111111100", xin_1 => "001000011110001001", pass => false),
  (xin_0 => "001000100010100110", xin_1 => "001011010000000110", pass => false),
  (xin_0 => "001010010010100110", xin_1 => "001011111110100110", pass => false),
  (xin_0 => "001001111110001000", xin_1 => "000110000110101111", pass => true),
  (xin_0 => "000100001100010011", xin_1 => "001000100011101100", pass => false),
  (xin_0 => "001000111110010100", xin_1 => "000011011010110011", pass => false),
  (xin_0 => "000111110001110111", xin_1 => "000010011010110011", pass => false),
  (xin_0 => "000011111010101000", xin_1 => "001000010110000100", pass => false),
  (xin_0 => "000111001010011010", xin_1 => "000100101100000111", pass => true),
  (xin_0 => "000100110001111010", xin_1 => "000101001000110101", pass => true),
  (xin_0 => "000111111110111110", xin_1 => "001011001011100000", pass => false),
  (xin_0 => "001000001101100001", xin_1 => "001010110110110100", pass => false),
  (xin_0 => "000011100010110010", xin_1 => "000010011001100000", pass => true),
  (xin_0 => "001011010011011101", xin_1 => "001001011111100010", pass => false),
  (xin_0 => "001001010110001110", xin_1 => "000001101101001001", pass => false),
  (xin_0 => "001100010111010000", xin_1 => "000111100001000011", pass => false),
  (xin_0 => "000110101011100100", xin_1 => "001011101101111101", pass => false),
  (xin_0 => "001000001110111001", xin_1 => "000110010011000111", pass => true),
  (xin_0 => "001101100000100110", xin_1 => "000101111000010111", pass => false),
  (xin_0 => "000101100010101000", xin_1 => "001000110110001100", pass => false),
  (xin_0 => "001010000001111000", xin_1 => "000100011100000011", pass => true),
  (xin_0 => "000011111011011011", xin_1 => "000101011111011100", pass => true),
  (xin_0 => "000011101000100010", xin_1 => "000101000111011100", pass => true),
  (xin_0 => "000100111110001110", xin_1 => "001000001100101100", pass => false),
  (xin_0 => "001110101100001010", xin_1 => "001010000110011011", pass => true),
  (xin_0 => "000011000100100111", xin_1 => "000001001100100110", pass => true),
  (xin_0 => "000110100001101000", xin_1 => "000010101011101101", pass => false),
  (xin_0 => "001000011101011101", xin_1 => "001001110011100011", pass => false),
  (xin_0 => "001100111000100101", xin_1 => "000011000000010100", pass => true),
  (xin_0 => "000110110110101101", xin_1 => "000001101110001100", pass => false),
  (xin_0 => "001011101000000011", xin_1 => "001001000011011011", pass => false),
  (xin_0 => "001101011000001111", xin_1 => "000000101111010011", pass => true),
  (xin_0 => "000100001001110001", xin_1 => "001000110000111011", pass => false),
  (xin_0 => "001010000100111110", xin_1 => "000101111110000000", pass => true),
  (xin_0 => "000110001000001011", xin_1 => "000101011001010111", pass => true),
  (xin_0 => "000111011101110001", xin_1 => "000010111110000010", pass => false),
  (xin_0 => "000111001010101011", xin_1 => "000011000111101110", pass => false),
  (xin_0 => "000011101011001000", xin_1 => "000101001100001001", pass => true),
  (xin_0 => "001001001011100101", xin_1 => "001011001011101010", pass => false),
  (xin_0 => "000011100001111000", xin_1 => "000011110110110010", pass => true),
  (xin_0 => "000110000001000011", xin_1 => "000001110001010100", pass => false),
  (xin_0 => "001001110001101011", xin_1 => "001101001111001101", pass => false),
  (xin_0 => "000110001100000001", xin_1 => "000010100110111000", pass => false),
  (xin_0 => "001011111101011010", xin_1 => "001000100110000111", pass => false),
  (xin_0 => "001000000110111010", xin_1 => "000010001101100001", pass => false),
  (xin_0 => "001100000000011101", xin_1 => "001001011110100110", pass => false),
  (xin_0 => "001100000010010100", xin_1 => "001000110010011100", pass => false),
  (xin_0 => "001011100101101111", xin_1 => "001000010000000001", pass => false),
  (xin_0 => "001001010101101111", xin_1 => "000101100010010101", pass => true),
  (xin_0 => "001101001011011100", xin_1 => "000001010100011100", pass => true),
  (xin_0 => "001100100111111110", xin_1 => "001000100101011001", pass => false),
  (xin_0 => "000111000010101110", xin_1 => "000010010111111001", pass => false),
  (xin_0 => "001100011011101100", xin_1 => "000111000110001011", pass => false),
  (xin_0 => "001100010111001001", xin_1 => "000110110110001110", pass => false),
  (xin_0 => "001010010111111100", xin_1 => "000110000101010010", pass => true),
  (xin_0 => "001001011011111011", xin_1 => "001000110111110111", pass => false),
  (xin_0 => "000110010011000010", xin_1 => "000011100110101110", pass => false),
  (xin_0 => "001000001111011010", xin_1 => "000011111110110100", pass => false),
  (xin_0 => "000111100011111011", xin_1 => "000110011000011100", pass => true),
  (xin_0 => "000111100111001001", xin_1 => "000110010011000011", pass => true),
  (xin_0 => "000111110100011010", xin_1 => "000100100100000111", pass => true),
  (xin_0 => "001011000011011011", xin_1 => "000011001110000000", pass => true),
  (xin_0 => "001100111001000111", xin_1 => "000101110111101110", pass => false),
  (xin_0 => "000101001001111101", xin_1 => "000101001001110001", pass => true),
  (xin_0 => "000101101011110111", xin_1 => "001000001101101111", pass => false),
  (xin_0 => "000011001010101110", xin_1 => "000110000010011011", pass => false),
  (xin_0 => "000110010000001111", xin_1 => "000011000111101010", pass => false),
  (xin_0 => "001011010111110000", xin_1 => "001001000010100011", pass => false),
  (xin_0 => "000111101001011110", xin_1 => "000011011001111101", pass => false),
  (xin_0 => "000110110000110001", xin_1 => "000100001010011111", pass => false),
  (xin_0 => "001011101001110010", xin_1 => "000111110000000101", pass => false),
  (xin_0 => "001000101011100101", xin_1 => "001011010100111101", pass => false),
  (xin_0 => "000100001101100010", xin_1 => "000000110001001001", pass => true),
  (xin_0 => "001101100000111110", xin_1 => "000101111100111001", pass => false),
  (xin_0 => "001010101001001110", xin_1 => "000101100101011000", pass => true),
  (xin_0 => "000100111011010100", xin_1 => "000010111001111101", pass => true),
  (xin_0 => "001100010001000001", xin_1 => "001000000100101001", pass => false),
  (xin_0 => "001010001000110110", xin_1 => "000001101001001000", pass => false),
  (xin_0 => "000111000000000110", xin_1 => "000100010101110110", pass => true),
  (xin_0 => "000100101010010111", xin_1 => "000010011111001010", pass => true),
  (xin_0 => "000111100010001111", xin_1 => "000010110001111001", pass => false),
  (xin_0 => "000111000111111001", xin_1 => "001010010101001111", pass => false),
  (xin_0 => "001001000001100000", xin_1 => "000100000010101110", pass => false),
  (xin_0 => "000110011010111001", xin_1 => "001001000001111011", pass => false),
  (xin_0 => "001010100010001001", xin_1 => "000101101110100000", pass => true),
  (xin_0 => "000100110010010000", xin_1 => "000100110011000011", pass => true),
  (xin_0 => "001000010001010001", xin_1 => "000010101010100101", pass => false),
  (xin_0 => "001101110001101111", xin_1 => "000110111101110111", pass => false),
  (xin_0 => "001011110001110001", xin_1 => "001000101011111001", pass => false),
  (xin_0 => "001001110110101100", xin_1 => "001011010100111000", pass => false),
  (xin_0 => "001010000001011001", xin_1 => "000111100001111011", pass => true),
  (xin_0 => "000110010011111110", xin_1 => "000100110000011111", pass => true),
  (xin_0 => "000101001100101010", xin_1 => "001000110111001101", pass => false),
  (xin_0 => "000101110001100100", xin_1 => "000010101011011110", pass => false),
  (xin_0 => "001000001011010001", xin_1 => "000010011010001000", pass => false),
  (xin_0 => "000110001001011101", xin_1 => "000011011101001110", pass => false),
  (xin_0 => "000101111100101001", xin_1 => "001001000100110011", pass => false),
  (xin_0 => "001001000100111010", xin_1 => "000010101001010010", pass => false),
  (xin_0 => "001000101010000101", xin_1 => "000101010010111110", pass => true),
  (xin_0 => "000111110000011111", xin_1 => "000110001001001110", pass => true),
  (xin_0 => "000110111100000011", xin_1 => "000011111111011001", pass => false),
  (xin_0 => "001001100010101101", xin_1 => "001000000110101001", pass => true),
  (xin_0 => "001100100010100000", xin_1 => "000111001010111100", pass => false),
  (xin_0 => "000111111100100101", xin_1 => "000001101011000001", pass => false),
  (xin_0 => "001000000001001001", xin_1 => "000101100101000010", pass => true),
  (xin_0 => "000101100010000010", xin_1 => "000011111011000010", pass => true),
  (xin_0 => "001001110000010011", xin_1 => "000101001111011111", pass => true),
  (xin_0 => "001011001010101000", xin_1 => "000011110010000110", pass => true),
  (xin_0 => "000010101110110110", xin_1 => "000011100111101101", pass => true),
  (xin_0 => "001010101010101101", xin_1 => "001001101111000000", pass => false),
  (xin_0 => "001000010100010110", xin_1 => "000101101000100101", pass => true),
  (xin_0 => "001010000100101100", xin_1 => "001011011100001010", pass => false),
  (xin_0 => "000101001011101001", xin_1 => "000010111100000110", pass => true),
  (xin_0 => "001011100101101100", xin_1 => "001000110110101100", pass => false),
  (xin_0 => "000111100111001001", xin_1 => "000010100101011101", pass => false),
  (xin_0 => "000100011101010000", xin_1 => "000011111101110110", pass => true),
  (xin_0 => "001110111011110001", xin_1 => "000011100000110000", pass => false),
  (xin_0 => "001011011101110110", xin_1 => "000010100111010101", pass => true),
  (xin_0 => "001001101000011111", xin_1 => "001001001000111111", pass => false),
  (xin_0 => "001101011011111000", xin_1 => "001001100101000011", pass => true),
  (xin_0 => "000011110010011001", xin_1 => "000101011101010101", pass => true),
  (xin_0 => "001011010101110101", xin_1 => "000111100110001101", pass => false),
  (xin_0 => "000110001101110100", xin_1 => "000001110111100000", pass => false),
  (xin_0 => "000110010011011111", xin_1 => "000111100001001011", pass => true),
  (xin_0 => "000110011010011100", xin_1 => "000010111100001011", pass => false),
  (xin_0 => "001001000111000110", xin_1 => "000001011001000011", pass => false),
  (xin_0 => "001110101101101011", xin_1 => "001001110100001111", pass => true),
  (xin_0 => "000100110101000010", xin_1 => "000100010110100100", pass => true),
  (xin_0 => "001010010011001001", xin_1 => "001000110010010111", pass => false),
  (xin_0 => "001101001010000011", xin_1 => "000110101111011001", pass => false),
  (xin_0 => "001010000010100111", xin_1 => "001010000110010010", pass => false),
  (xin_0 => "001011111000111111", xin_1 => "000111000000100110", pass => false),
  (xin_0 => "001000001011001100", xin_1 => "001011000101110101", pass => false),
  (xin_0 => "001101000001000101", xin_1 => "000010110011001011", pass => true),
  (xin_0 => "001000101011011001", xin_1 => "000011101110111001", pass => false),
  (xin_0 => "000110100011100110", xin_1 => "001001111110000001", pass => false),
  (xin_0 => "001010111001010010", xin_1 => "001001101110101010", pass => false),
  (xin_0 => "001001001111001100", xin_1 => "000111101000111100", pass => true),
  (xin_0 => "000110110000100001", xin_1 => "000010100011101001", pass => false),
  (xin_0 => "000100110111000111", xin_1 => "000101001001000010", pass => true),
  (xin_0 => "000101000110101000", xin_1 => "000100011101100100", pass => true),
  (xin_0 => "000011000010000110", xin_1 => "000100011101000011", pass => true),
  (xin_0 => "001010101101000101", xin_1 => "000111010111010110", pass => false),
  (xin_0 => "001001000111110110", xin_1 => "000101000101000101", pass => true),
  (xin_0 => "000101110001101101", xin_1 => "000110101010101111", pass => true),
  (xin_0 => "001100010011011111", xin_1 => "000010010010000001", pass => true),
  (xin_0 => "001000110010001100", xin_1 => "000010101110100000", pass => false),
  (xin_0 => "000100100100111110", xin_1 => "000111011001001111", pass => false),
  (xin_0 => "000110110100110011", xin_1 => "000010100111010101", pass => false),
  (xin_0 => "000110001000001001", xin_1 => "001000011011100110", pass => false),
  (xin_0 => "001111100110001110", xin_1 => "001010001110110001", pass => true),
  (xin_0 => "001001111110110100", xin_1 => "000101100011010100", pass => true),
  (xin_0 => "000100101110010111", xin_1 => "000101111001100010", pass => true),
  (xin_0 => "001111011000110010", xin_1 => "001010001110010000", pass => true),
  (xin_0 => "001100101000001001", xin_1 => "000101101111101011", pass => false),
  (xin_0 => "000100100111111001", xin_1 => "000100101101101011", pass => true),
  (xin_0 => "001100000110110011", xin_1 => "000101000011111101", pass => true),
  (xin_0 => "001011110011011000", xin_1 => "001000000101010111", pass => false),
  (xin_0 => "001000000100010000", xin_1 => "001101001001011000", pass => false),
  (xin_0 => "001011101010111101", xin_1 => "000101011100111010", pass => true),
  (xin_0 => "001100111101011011", xin_1 => "000011001000110101", pass => true),
  (xin_0 => "001000001000001110", xin_1 => "001100010000011100", pass => false),
  (xin_0 => "001100011101110110", xin_1 => "000010011110000001", pass => true),
  (xin_0 => "001000010101110110", xin_1 => "000100010010101100", pass => false),
  (xin_0 => "001001000000010001", xin_1 => "000110100000101100", pass => true),
  (xin_0 => "000100011100111000", xin_1 => "001000000000111011", pass => false),
  (xin_0 => "001000000011100011", xin_1 => "000010011000000011", pass => false),
  (xin_0 => "001000110000010110", xin_1 => "000101000000000100", pass => true),
  (xin_0 => "000100010110010101", xin_1 => "001000100010111111", pass => false),
  (xin_0 => "000011011100001010", xin_1 => "001000110101001010", pass => false),
  (xin_0 => "000111111001011110", xin_1 => "000001111101110111", pass => false),
  (xin_0 => "001000001001111000", xin_1 => "001001011011000110", pass => false),
  (xin_0 => "000110010110010001", xin_1 => "000110011010101001", pass => true),
  (xin_0 => "000101100111000110", xin_1 => "000100001110011100", pass => true),
  (xin_0 => "001001110111101110", xin_1 => "000110001010000010", pass => true),
  (xin_0 => "000111111001000110", xin_1 => "000011100011000011", pass => false),
  (xin_0 => "001101110010100001", xin_1 => "000110011111101000", pass => false),
  (xin_0 => "001001011000110110", xin_1 => "000101011100110001", pass => true),
  (xin_0 => "000110011000001001", xin_1 => "000011100010100100", pass => false),
  (xin_0 => "001101000110100100", xin_1 => "000111101100101000", pass => false),
  (xin_0 => "001000010111110000", xin_1 => "000110011100101100", pass => true),
  (xin_0 => "000101110100000011", xin_1 => "001001110101100010", pass => false),
  (xin_0 => "001011111111111111", xin_1 => "000100000001110111", pass => true),
  (xin_0 => "000101011000011100", xin_1 => "001000111011101000", pass => false),
  (xin_0 => "001010100011100101", xin_1 => "001010111010010101", pass => false),
  (xin_0 => "000110111000100001", xin_1 => "000010000110011010", pass => false),
  (xin_0 => "001011110101101110", xin_1 => "000001000100001100", pass => true),
  (xin_0 => "001000101110010110", xin_1 => "000010000010101111", pass => false),
  (xin_0 => "001011110001110110", xin_1 => "001010101101110100", pass => false),
  (xin_0 => "000101011101101010", xin_1 => "000010100110110101", pass => false),
  (xin_0 => "000011110011101000", xin_1 => "000010111101011100", pass => true),
  (xin_0 => "000100011010110010", xin_1 => "000101101101001000", pass => true),
  (xin_0 => "001101100011100110", xin_1 => "000101111011110101", pass => false),
  (xin_0 => "000100101000001000", xin_1 => "000110001101111011", pass => true),
  (xin_0 => "000111110100111100", xin_1 => "000010001110101011", pass => false),
  (xin_0 => "000011010000000010", xin_1 => "000101011001110101", pass => true),
  (xin_0 => "000111010101110110", xin_1 => "000100101100010111", pass => true),
  (xin_0 => "000100111111101111", xin_1 => "001000001011111101", pass => false),
  (xin_0 => "000111100111010000", xin_1 => "000101101010001011", pass => true),
  (xin_0 => "001001111001001111", xin_1 => "000101110000110011", pass => true),
  (xin_0 => "001001001100001110", xin_1 => "000101000001000110", pass => true),
  (xin_0 => "000111100010110010", xin_1 => "000001010011100011", pass => false),
  (xin_0 => "000101111001011100", xin_1 => "001000011010100101", pass => false),
  (xin_0 => "000110111000101010", xin_1 => "000101101111010001", pass => true),
  (xin_0 => "001101011100001011", xin_1 => "000110001000101000", pass => false),
  (xin_0 => "001011100110100000", xin_1 => "000111000001000101", pass => false),
  (xin_0 => "000011010000011111", xin_1 => "000100001011100000", pass => true),
  (xin_0 => "001000011110110001", xin_1 => "000011111010111101", pass => false),
  (xin_0 => "000110101100010111", xin_1 => "000010000100010101", pass => false),
  (xin_0 => "001000011100100001", xin_1 => "000011011101101110", pass => false),
  (xin_0 => "001011110000110011", xin_1 => "001001101101110000", pass => false),
  (xin_0 => "001011010000010100", xin_1 => "001001010010101000", pass => false),
  (xin_0 => "000110011111000100", xin_1 => "001010001110111000", pass => false),
  (xin_0 => "001100100010000000", xin_1 => "001100111000110000", pass => false),
  (xin_0 => "001011011101100101", xin_1 => "001001101011011001", pass => false),
  (xin_0 => "000110000110110011", xin_1 => "000010111100111100", pass => false),
  (xin_0 => "001010100011011111", xin_1 => "000101101101000100", pass => true),
  (xin_0 => "001000110000101110", xin_1 => "000100110001010111", pass => true),
  (xin_0 => "001101100011110010", xin_1 => "001011011100100100", pass => true),
  (xin_0 => "001001011011100111", xin_1 => "000100111111110110", pass => true),
  (xin_0 => "000100100010111100", xin_1 => "000100001110101000", pass => true),
  (xin_0 => "001101101001000000", xin_1 => "000010101101100000", pass => true),
  (xin_0 => "000110101000011010", xin_1 => "001011101000110111", pass => false),
  (xin_0 => "000110010110001111", xin_1 => "000010000010101001", pass => false),
  (xin_0 => "001001111000010110", xin_1 => "000011001100011011", pass => false),
  (xin_0 => "001101101101111010", xin_1 => "000110110000011110", pass => false),
  (xin_0 => "000110001010101101", xin_1 => "001001010001010110", pass => false),
  (xin_0 => "000010011011110001", xin_1 => "000110101111000011", pass => false),
  (xin_0 => "001100011010011001", xin_1 => "000111000110110100", pass => false),
  (xin_0 => "001011101010011010", xin_1 => "000111111010101111", pass => false),
  (xin_0 => "001101111101111001", xin_1 => "001011010110000011", pass => true),
  (xin_0 => "001010000011010111", xin_1 => "001011100001110101", pass => false),
  (xin_0 => "001100101011101010", xin_1 => "000111110100101001", pass => false),
  (xin_0 => "000111001110000100", xin_1 => "000010000111101001", pass => false),
  (xin_0 => "000111000011110010", xin_1 => "000011001000000111", pass => false),
  (xin_0 => "000101010111000100", xin_1 => "001001010001101101", pass => false),
  (xin_0 => "000111111111110110", xin_1 => "000110011110101100", pass => true),
  (xin_0 => "001001000111011010", xin_1 => "000100110001011010", pass => true),
  (xin_0 => "001001110000111110", xin_1 => "000111100010000101", pass => true),
  (xin_0 => "001001000000010000", xin_1 => "001010101011111101", pass => false),
  (xin_0 => "000011110101111111", xin_1 => "000010101011001100", pass => true),
  (xin_0 => "001101011101010111", xin_1 => "000100110011111001", pass => false),
  (xin_0 => "001010001111011101", xin_1 => "000010000001100010", pass => false),
  (xin_0 => "000111100000100011", xin_1 => "000011111001100001", pass => false),
  (xin_0 => "000111010011010000", xin_1 => "000111110000001011", pass => true),
  (xin_0 => "000111000010100100", xin_1 => "000110000000110010", pass => true),
  (xin_0 => "001000100011011000", xin_1 => "000010000100000100", pass => false),
  (xin_0 => "001010011001010011", xin_1 => "000011000111011100", pass => false),
  (xin_0 => "001100000110011000", xin_1 => "001000000011011001", pass => false),
  (xin_0 => "001100011111010011", xin_1 => "000110001011001101", pass => false),
  (xin_0 => "000100110011011100", xin_1 => "000011000111011100", pass => true),
  (xin_0 => "000111110100110110", xin_1 => "000010100101010001", pass => false),
  (xin_0 => "000111101011100010", xin_1 => "000111001110111011", pass => true),
  (xin_0 => "001101111011100100", xin_1 => "000110010100001110", pass => false),
  (xin_0 => "001000101001110111", xin_1 => "000110010101101111", pass => true),
  (xin_0 => "001000000101110000", xin_1 => "000010011001100010", pass => false),
  (xin_0 => "001000010001011000", xin_1 => "000010100001111100", pass => false),
  (xin_0 => "001101001111011011", xin_1 => "001011101000000111", pass => true),
  (xin_0 => "001101100101110111", xin_1 => "000010000101011110", pass => true),
  (xin_0 => "001101110111101111", xin_1 => "000100101111011001", pass => false),
  (xin_0 => "001101001001011011", xin_1 => "000111011100000001", pass => false),
  (xin_0 => "000111000000010001", xin_1 => "000111001011011110", pass => true),
  (xin_0 => "001000100000100111", xin_1 => "000010100100111110", pass => false),
  (xin_0 => "001100011111101100", xin_1 => "000111001101101111", pass => false),
  (xin_0 => "000101111011101101", xin_1 => "001010000100101111", pass => false),
  (xin_0 => "000100111110010001", xin_1 => "001000101011101100", pass => false),
  (xin_0 => "001100111100101111", xin_1 => "001000010110010100", pass => false),
  (xin_0 => "001101010111110100", xin_1 => "000111010011110001", pass => false),
  (xin_0 => "000101001001110110", xin_1 => "000110001111111110", pass => true),
  (xin_0 => "001111101100100010", xin_1 => "001001111001001011", pass => true),
  (xin_0 => "000100010101111101", xin_1 => "000011001111111001", pass => true),
  (xin_0 => "001001011001101100", xin_1 => "000110010101110100", pass => true),
  (xin_0 => "000111100000001011", xin_1 => "000001110111011001", pass => false),
  (xin_0 => "000110000000111110", xin_1 => "000010000101101111", pass => false),
  (xin_0 => "001011001010011000", xin_1 => "000101001101101010", pass => true),
  (xin_0 => "000110111010110010", xin_1 => "000010100101001000", pass => false),
  (xin_0 => "001100011110100110", xin_1 => "000001110010101111", pass => true),
  (xin_0 => "001010000111110001", xin_1 => "000110010100010110", pass => true),
  (xin_0 => "000011011101011100", xin_1 => "000010111000011100", pass => true),
  (xin_0 => "000111001111100110", xin_1 => "000101001110101011", pass => true),
  (xin_0 => "001000010110100100", xin_1 => "000011111101100111", pass => false),
  (xin_0 => "001100101000100010", xin_1 => "001000000001000111", pass => false),
  (xin_0 => "001001001111111100", xin_1 => "000010000101100000", pass => false),
  (xin_0 => "001011001101111111", xin_1 => "000101110011100000", pass => true),
  (xin_0 => "001101001100010111", xin_1 => "000110000101100001", pass => false),
  (xin_0 => "000110111000011100", xin_1 => "000110011111010001", pass => true),
  (xin_0 => "001010100001000101", xin_1 => "000010011001001101", pass => false),
  (xin_0 => "001011011001111100", xin_1 => "001011111010000100", pass => false),
  (xin_0 => "000011111101001010", xin_1 => "000100111110101101", pass => true),
  (xin_0 => "000100111011011001", xin_1 => "000010000111000110", pass => true),
  (xin_0 => "000111101001101101", xin_1 => "001001011001000110", pass => false),
  (xin_0 => "001001100011100010", xin_1 => "000100111011011010", pass => true),
  (xin_0 => "001001000000011000", xin_1 => "001011010100101101", pass => false),
  (xin_0 => "000110110110110010", xin_1 => "000010011001101101", pass => false),
  (xin_0 => "001010110010111101", xin_1 => "001000100001100100", pass => false),
  (xin_0 => "001011000011010011", xin_1 => "001001001110111011", pass => false),
  (xin_0 => "000101000111101001", xin_1 => "001000111111000001", pass => false),
  (xin_0 => "001010010110100010", xin_1 => "000010011111010100", pass => false),
  (xin_0 => "000111011101101111", xin_1 => "000010100011000001", pass => false),
  (xin_0 => "001010110011100110", xin_1 => "001001110111011000", pass => false),
  (xin_0 => "001001001010011100", xin_1 => "001000000010100100", pass => true),
  (xin_0 => "000111100100010110", xin_1 => "000011110011100111", pass => false),
  (xin_0 => "001001101101100100", xin_1 => "000100100101111011", pass => true),
  (xin_0 => "001001110111000111", xin_1 => "000010111111000000", pass => false),
  (xin_0 => "001100100000101100", xin_1 => "000101111101100011", pass => false),
  (xin_0 => "001001010111100000", xin_1 => "000011110101101110", pass => false),
  (xin_0 => "000111011000011101", xin_1 => "001001000001010000", pass => false),
  (xin_0 => "000110010100001000", xin_1 => "000011011101111101", pass => false),
  (xin_0 => "001000000110100010", xin_1 => "000001100010100111", pass => false),
  (xin_0 => "001001011000110000", xin_1 => "001010001011010100", pass => false),
  (xin_0 => "000110111011100000", xin_1 => "000010011000110111", pass => false),
  (xin_0 => "001000110010001010", xin_1 => "000111110111101100", pass => true),
  (xin_0 => "001000000000010000", xin_1 => "000110111011100111", pass => true),
  (xin_0 => "000101100001101011", xin_1 => "000100101001000010", pass => true),
  (xin_0 => "000111111100101111", xin_1 => "000010101110101101", pass => false),
  (xin_0 => "001100001000101010", xin_1 => "000111110001010100", pass => false),
  (xin_0 => "001000110010001111", xin_1 => "000011011110101101", pass => false),
  (xin_0 => "000111000100000001", xin_1 => "001001101100010101", pass => false),
  (xin_0 => "000010111101010001", xin_1 => "000100101001001001", pass => true),
  (xin_0 => "000101110111110011", xin_1 => "000111101111001000", pass => true),
  (xin_0 => "001011001100110001", xin_1 => "000110010001111001", pass => true),
  (xin_0 => "001101011001010001", xin_1 => "000111010110001001", pass => false),
  (xin_0 => "001101100000110010", xin_1 => "000110101111110110", pass => false),
  (xin_0 => "001100011000100101", xin_1 => "000011011100001110", pass => true),
  (xin_0 => "000101001100100100", xin_1 => "001001110000010010", pass => false),
  (xin_0 => "001000010011110011", xin_1 => "000110101100111101", pass => true),
  (xin_0 => "000110100001010111", xin_1 => "000110100100000111", pass => true),
  (xin_0 => "000101110110000010", xin_1 => "000110001011010000", pass => true),
  (xin_0 => "001000001011010000", xin_1 => "000001100110110101", pass => false),
  (xin_0 => "000111011111001100", xin_1 => "000010111010101100", pass => false),
  (xin_0 => "001010001010111110", xin_1 => "001100100111001000", pass => false),
  (xin_0 => "001001010100111100", xin_1 => "001010110110010011", pass => false),
  (xin_0 => "001000000110110101", xin_1 => "000101100010111110", pass => true),
  (xin_0 => "000110111110111000", xin_1 => "001011010110000100", pass => false),
  (xin_0 => "001001111110111001", xin_1 => "001100100010101111", pass => false),
  (xin_0 => "000111001011011111", xin_1 => "000001111010110010", pass => false),
  (xin_0 => "010000000010110111", xin_1 => "001010000001110100", pass => true),
  (xin_0 => "001001101000001100", xin_1 => "000010010011010000", pass => false),
  (xin_0 => "001011100100111001", xin_1 => "000100100011010101", pass => true),
  (xin_0 => "001000010110110111", xin_1 => "000110001010100010", pass => true),
  (xin_0 => "001011100001111000", xin_1 => "000100100000100000", pass => true),
  (xin_0 => "001000110110101010", xin_1 => "000110101010101100", pass => true),
  (xin_0 => "001010000100100100", xin_1 => "000011001100100110", pass => false),
  (xin_0 => "001010001101101001", xin_1 => "000111011011110011", pass => true),
  (xin_0 => "001001010111011111", xin_1 => "000001011111011111", pass => false),
  (xin_0 => "001011010100100101", xin_1 => "000011010111011101", pass => true),
  (xin_0 => "000100001111111111", xin_1 => "000111101001101101", pass => false),
  (xin_0 => "001011110101100110", xin_1 => "000001010000110010", pass => true),
  (xin_0 => "001010011011111101", xin_1 => "000010001010100011", pass => false),
  (xin_0 => "001000010101100001", xin_1 => "000111000000111011", pass => true),
  (xin_0 => "000111101010110001", xin_1 => "001001010101000011", pass => false),
  (xin_0 => "000111011011111010", xin_1 => "000010111011000111", pass => false),
  (xin_0 => "000110010111100001", xin_1 => "001001010100001111", pass => false),
  (xin_0 => "001011011111000101", xin_1 => "001011101010110011", pass => false),
  (xin_0 => "001010100110011101", xin_1 => "000100100101110110", pass => true),
  (xin_0 => "001011011111110011", xin_1 => "000010000001111111", pass => true),
  (xin_0 => "001010000010011111", xin_1 => "001001111111101010", pass => false),
  (xin_0 => "001010011111111110", xin_1 => "000011111010000101", pass => true),
  (xin_0 => "001000110000011000", xin_1 => "000010011110000010", pass => false),
  (xin_0 => "001101000110111111", xin_1 => "000110101011001010", pass => false),
  (xin_0 => "000010111100000011", xin_1 => "000000110011101001", pass => true),
  (xin_0 => "001001001011100111", xin_1 => "000101111011001001", pass => true),
  (xin_0 => "001011111111110111", xin_1 => "000100110011110010", pass => true),
  (xin_0 => "001001000100101010", xin_1 => "000111010001101101", pass => true),
  (xin_0 => "001100101000110101", xin_1 => "000111101110111110", pass => false),
  (xin_0 => "000111000101000111", xin_1 => "001001100000011100", pass => false),
  (xin_0 => "000110100001010000", xin_1 => "000010101100010111", pass => false),
  (xin_0 => "001001100100011010", xin_1 => "001011101110000101", pass => false),
  (xin_0 => "001010100001011000", xin_1 => "001010100000001010", pass => false),
  (xin_0 => "000101001010001001", xin_1 => "000010101101100000", pass => true),
  (xin_0 => "001010111110011011", xin_1 => "001000100111000001", pass => false),
  (xin_0 => "000110111100101100", xin_1 => "001000100010001011", pass => true),
  (xin_0 => "000111010101001010", xin_1 => "001001011101000010", pass => false),
  (xin_0 => "001010001100011110", xin_1 => "000100101110011110", pass => true),
  (xin_0 => "000100001111111111", xin_1 => "001001010101110111", pass => false),
  (xin_0 => "000100101011101110", xin_1 => "000101100101001111", pass => true),
  (xin_0 => "000110110001110010", xin_1 => "000010000011111011", pass => false),
  (xin_0 => "001001110011110100", xin_1 => "001010110101001010", pass => false),
  (xin_0 => "000111010000110100", xin_1 => "000011111110000000", pass => false),
  (xin_0 => "001010001010011110", xin_1 => "000010110011110101", pass => false),
  (xin_0 => "000011111111000001", xin_1 => "000100001111011110", pass => true),
  (xin_0 => "000111111110101110", xin_1 => "000110000100011000", pass => true),
  (xin_0 => "000111000111101101", xin_1 => "000111000000100010", pass => true),
  (xin_0 => "000110011001011010", xin_1 => "000100000001010010", pass => false),
  (xin_0 => "001000100000111111", xin_1 => "001011010001111111", pass => false),
  (xin_0 => "000110111110111111", xin_1 => "000010111101110110", pass => false),
  (xin_0 => "001010110011001110", xin_1 => "001001100110110010", pass => false),
  (xin_0 => "001100100111111001", xin_1 => "000111101110100011", pass => false),
  (xin_0 => "001110111101001101", xin_1 => "001010011000001111", pass => true),
  (xin_0 => "001101110010011001", xin_1 => "000000110111000000", pass => true),
  (xin_0 => "001010010011101111", xin_1 => "001001001110010100", pass => false),
  (xin_0 => "000110011010011010", xin_1 => "000101000000011101", pass => true),
  (xin_0 => "001001011101011111", xin_1 => "001000001101010100", pass => true),
  (xin_0 => "000111010110111011", xin_1 => "000110111100011111", pass => true),
  (xin_0 => "001100010011001111", xin_1 => "001000000010110110", pass => false),
  (xin_0 => "000101010000101111", xin_1 => "000100001000101110", pass => true),
  (xin_0 => "000111000100010011", xin_1 => "001001101001010110", pass => false),
  (xin_0 => "001001010100010110", xin_1 => "001000101101110111", pass => false),
  (xin_0 => "000101101110111111", xin_1 => "000111001010100101", pass => true),
  (xin_0 => "001101010111000010", xin_1 => "000110000001110111", pass => false),
  (xin_0 => "000111110110010010", xin_1 => "000010111011110001", pass => false),
  (xin_0 => "000111000111100101", xin_1 => "000010101000110100", pass => false),
  (xin_0 => "000101011101000100", xin_1 => "000011101000010111", pass => true),
  (xin_0 => "001011111111110010", xin_1 => "000100001111001100", pass => true),
  (xin_0 => "001011100100100001", xin_1 => "000101001100101001", pass => true),
  (xin_0 => "000111000000110101", xin_1 => "001001111011101001", pass => false),
  (xin_0 => "000110100010010010", xin_1 => "000101011100010110", pass => true),
  (xin_0 => "001100001011011000", xin_1 => "000111111101010111", pass => false),
  (xin_0 => "000110011011111001", xin_1 => "000110000110111011", pass => true),
  (xin_0 => "000100011101111100", xin_1 => "001001011010110011", pass => false),
  (xin_0 => "001110110101111011", xin_1 => "001010001111110100", pass => true),
  (xin_0 => "001001011101101111", xin_1 => "000010111110001000", pass => false),
  (xin_0 => "001010001110101010", xin_1 => "000110111110011110", pass => true),
  (xin_0 => "000100101000000001", xin_1 => "000111011111010011", pass => false),
  (xin_0 => "001000011000100010", xin_1 => "000111111000011011", pass => true),
  (xin_0 => "000101010101001111", xin_1 => "000010110001101110", pass => true),
  (xin_0 => "001000100110111010", xin_1 => "000011101010101101", pass => false),
  (xin_0 => "001100010100000101", xin_1 => "001000010111010000", pass => false),
  (xin_0 => "000101010101111011", xin_1 => "000110100010110001", pass => true),
  (xin_0 => "001111011010011000", xin_1 => "001000111100100101", pass => true),
  (xin_0 => "001010000100111100", xin_1 => "001011001100111100", pass => false),
  (xin_0 => "000011101111010000", xin_1 => "001000010010001000", pass => false),
  (xin_0 => "001010101010110011", xin_1 => "000110111100001111", pass => true),
  (xin_0 => "001001010011100110", xin_1 => "000110000110100110", pass => true),
  (xin_0 => "000011111011100111", xin_1 => "000010010001111000", pass => true),
  (xin_0 => "001100000100100010", xin_1 => "001000110001110000", pass => false),
  (xin_0 => "001011100100001001", xin_1 => "000011010101010011", pass => true),
  (xin_0 => "000110001100101000", xin_1 => "000010001011101110", pass => false),
  (xin_0 => "001001100000011101", xin_1 => "001100000111110011", pass => false),
  (xin_0 => "001010010000011110", xin_1 => "000101111010011000", pass => true),
  (xin_0 => "000011111111101011", xin_1 => "000101010000100100", pass => true),
  (xin_0 => "000111111111110011", xin_1 => "000111001001001001", pass => true),
  (xin_0 => "000110110011000010", xin_1 => "000100111101110011", pass => true),
  (xin_0 => "001001010100001100", xin_1 => "000010011101011000", pass => false),
  (xin_0 => "000111110110010111", xin_1 => "001010100000101001", pass => false),
  (xin_0 => "000100100010001111", xin_1 => "000110111110011101", pass => true),
  (xin_0 => "000111100011100111", xin_1 => "000110100000001001", pass => true),
  (xin_0 => "001100000111110100", xin_1 => "000100100101111100", pass => true),
  (xin_0 => "001100010010011011", xin_1 => "000001000110000010", pass => true),
  (xin_0 => "001011111110111100", xin_1 => "000110111001001010", pass => false),
  (xin_0 => "001010110100000001", xin_1 => "001000111111011011", pass => false),
  (xin_0 => "001011000111000111", xin_1 => "001000010011000111", pass => false),
  (xin_0 => "000110001011101100", xin_1 => "001001100110111100", pass => false),
  (xin_0 => "000011001110110111", xin_1 => "000001000000111001", pass => true),
  (xin_0 => "000111100110001001", xin_1 => "000010101011000001", pass => false),
  (xin_0 => "000101000111001011", xin_1 => "000110010110010011", pass => true),
  (xin_0 => "001110000111011111", xin_1 => "001010010101110000", pass => true),
  (xin_0 => "000111100110001101", xin_1 => "000110111110001101", pass => true),
  (xin_0 => "001001011100101001", xin_1 => "000011100010001011", pass => false),
  (xin_0 => "001100100010100100", xin_1 => "000110001111000001", pass => false),
  (xin_0 => "001000100011101001", xin_1 => "000010101100001011", pass => false),
  (xin_0 => "001010011001010011", xin_1 => "000111111100111010", pass => false),
  (xin_0 => "001001100000110110", xin_1 => "001011011101001101", pass => false),
  (xin_0 => "001100111110101111", xin_1 => "000110101100110010", pass => false),
  (xin_0 => "000011101010110001", xin_1 => "000011011111110000", pass => true),
  (xin_0 => "001101011110011010", xin_1 => "000101101100001001", pass => false),
  (xin_0 => "001010011000100101", xin_1 => "000011001001010000", pass => false),
  (xin_0 => "001001010110011011", xin_1 => "001011010110110000", pass => false),
  (xin_0 => "001011111100100100", xin_1 => "000110010101000000", pass => false),
  (xin_0 => "000101101100001111", xin_1 => "000110110100001101", pass => true),
  (xin_0 => "000101000100011100", xin_1 => "001000001000010111", pass => false),
  (xin_0 => "001001001101001000", xin_1 => "000010010110001000", pass => false),
  (xin_0 => "001000111110111101", xin_1 => "000010011001001011", pass => false),
  (xin_0 => "001111000001000010", xin_1 => "001001100100101010", pass => true),
  (xin_0 => "000101100000101101", xin_1 => "000010001110001010", pass => false),
  (xin_0 => "000111111110011100", xin_1 => "001010101111010110", pass => false),
  (xin_0 => "000110110000010001", xin_1 => "000111010101110011", pass => true),
  (xin_0 => "001001100001011010", xin_1 => "001001100000100011", pass => false),
  (xin_0 => "001010100011010111", xin_1 => "000101100111110110", pass => true),
  (xin_0 => "001011110010111010", xin_1 => "000110100000011110", pass => false),
  (xin_0 => "001010101011011011", xin_1 => "000111100001111101", pass => false),
  (xin_0 => "000101010111010001", xin_1 => "000011011011110000", pass => true),
  (xin_0 => "000100101000000101", xin_1 => "001000101001011111", pass => false),
  (xin_0 => "001011100110010100", xin_1 => "000001011000001101", pass => true),
  (xin_0 => "000110110100010000", xin_1 => "000110000001011001", pass => true),
  (xin_0 => "000111111000011000", xin_1 => "001010101110001100", pass => false),
  (xin_0 => "001100101011100011", xin_1 => "000001111000011001", pass => true),
  (xin_0 => "000111101001010110", xin_1 => "001011011100100011", pass => false),
  (xin_0 => "001001000111000111", xin_1 => "000010001110101010", pass => false),
  (xin_0 => "001000010010001001", xin_1 => "000011111100101100", pass => false),
  (xin_0 => "001110100010010010", xin_1 => "000011101010101100", pass => false),
  (xin_0 => "001001110110010100", xin_1 => "000011000101100101", pass => false),
  (xin_0 => "001010100111000100", xin_1 => "000010011100111110", pass => false),
  (xin_0 => "001011100110111010", xin_1 => "000110001001100110", pass => true),
  (xin_0 => "000100111000111011", xin_1 => "000101000011011010", pass => true),
  (xin_0 => "001100101111100100", xin_1 => "000110101111100101", pass => false),
  (xin_0 => "000111100000011001", xin_1 => "000010001111010110", pass => false),
  (xin_0 => "001000011011101010", xin_1 => "001000000010010001", pass => true),
  (xin_0 => "001001100010001011", xin_1 => "000100011000000110", pass => true),
  (xin_0 => "001001011111111000", xin_1 => "001001000000011000", pass => false),
  (xin_0 => "000101110100011010", xin_1 => "001000111011101000", pass => false),
  (xin_0 => "000110110001111011", xin_1 => "000011100011001100", pass => false),
  (xin_0 => "001010100101011101", xin_1 => "000110101001001000", pass => true),
  (xin_0 => "001110000111110001", xin_1 => "000100101011101100", pass => false),
  (xin_0 => "001010010111010100", xin_1 => "001010010001111110", pass => false),
  (xin_0 => "001000001100011101", xin_1 => "001010000111110101", pass => false),
  (xin_0 => "000111001111000011", xin_1 => "001010000111011111", pass => false),
  (xin_0 => "001010100100011000", xin_1 => "000101011101000010", pass => true),
  (xin_0 => "001000100010110111", xin_1 => "000101110111011111", pass => true),
  (xin_0 => "000101111101100100", xin_1 => "000110101100010011", pass => true),
  (xin_0 => "001010000110111100", xin_1 => "000001101111001101", pass => false),
  (xin_0 => "001111101110111101", xin_1 => "000010011010011111", pass => false),
  (xin_0 => "001011011010100110", xin_1 => "001000011011101101", pass => false),
  (xin_0 => "001111011110011101", xin_1 => "001001111001011010", pass => true),
  (xin_0 => "001101111010000101", xin_1 => "000110000110000000", pass => false),
  (xin_0 => "001011010111100000", xin_1 => "000101011101000100", pass => true),
  (xin_0 => "000011011101110000", xin_1 => "000011110011001000", pass => true),
  (xin_0 => "001100000110111111", xin_1 => "000001011001111111", pass => true),
  (xin_0 => "000110111111111100", xin_1 => "001000110010010011", pass => false),
  (xin_0 => "000111101101100011", xin_1 => "000100101011100100", pass => true),
  (xin_0 => "001010110100110001", xin_1 => "001000100101111101", pass => false),
  (xin_0 => "000110111110111010", xin_1 => "000111001011101010", pass => true),
  (xin_0 => "000111011010010100", xin_1 => "000101101011110011", pass => true),
  (xin_0 => "001000001010001010", xin_1 => "000011001101111110", pass => false),
  (xin_0 => "000111100010111000", xin_1 => "000011100001111101", pass => false),
  (xin_0 => "001011101010000101", xin_1 => "000101011000101011", pass => true),
  (xin_0 => "001000110100111110", xin_1 => "001000000100010000", pass => true),
  (xin_0 => "000111101000100000", xin_1 => "001010111011110011", pass => false),
  (xin_0 => "001100011101111101", xin_1 => "000110010000001011", pass => false),
  (xin_0 => "001000101001011100", xin_1 => "000111111001111011", pass => true),
  (xin_0 => "001011111111100000", xin_1 => "001000100100000001", pass => false),
  (xin_0 => "001011010101000011", xin_1 => "001011110011100011", pass => false),
  (xin_0 => "000011100111010111", xin_1 => "000010011111011000", pass => true),
  (xin_0 => "000111110100100001", xin_1 => "000110110001110101", pass => true),
  (xin_0 => "000110000000110101", xin_1 => "000001001101101011", pass => false),
  (xin_0 => "000100111000110110", xin_1 => "000101111001110010", pass => true),
  (xin_0 => "000101110101111111", xin_1 => "000100100011001000", pass => true),
  (xin_0 => "001010110111001000", xin_1 => "001010001000000001", pass => false),
  (xin_0 => "000100001010101111", xin_1 => "000100000000011010", pass => true),
  (xin_0 => "001011101001011010", xin_1 => "001000001100111101", pass => false),
  (xin_0 => "001000010100100011", xin_1 => "000011100011000000", pass => false),
  (xin_0 => "001100110111100110", xin_1 => "000101000011010111", pass => true),
  (xin_0 => "001011101110001010", xin_1 => "000101100001111001", pass => true),
  (xin_0 => "000101001110110101", xin_1 => "000111111011010111", pass => false),
  (xin_0 => "001110101010110000", xin_1 => "001010100001100011", pass => true),
  (xin_0 => "001010100010001110", xin_1 => "000101101000100010", pass => true),
  (xin_0 => "000011110010011111", xin_1 => "000100011111011000", pass => true),
  (xin_0 => "001100011111110110", xin_1 => "001000110000111001", pass => false),
  (xin_0 => "001110011001100000", xin_1 => "000110100101000101", pass => false),
  (xin_0 => "000111000101011100", xin_1 => "000101100000010000", pass => true),
  (xin_0 => "001001110010100111", xin_1 => "001000000010111011", pass => true),
  (xin_0 => "001000110100110010", xin_1 => "000101001101011100", pass => true),
  (xin_0 => "001001000110101111", xin_1 => "000011101000101011", pass => false),
  (xin_0 => "000111001111100010", xin_1 => "000011000011111110", pass => false),
  (xin_0 => "001000010100001100", xin_1 => "000010110101001010", pass => false),
  (xin_0 => "001001111110001100", xin_1 => "000001111011010001", pass => false),
  (xin_0 => "001011101001000010", xin_1 => "000101111010110001", pass => true),
  (xin_0 => "001010011110001111", xin_1 => "000100010000011111", pass => true),
  (xin_0 => "001010001010000000", xin_1 => "001011101100010001", pass => false),
  (xin_0 => "001100000111111000", xin_1 => "000010000011011101", pass => true),
  (xin_0 => "000100111110111001", xin_1 => "000110101011101111", pass => true),
  (xin_0 => "000101001100001111", xin_1 => "000111111110110111", pass => false),
  (xin_0 => "001010011110000000", xin_1 => "000010000001011010", pass => false),
  (xin_0 => "001100000100110100", xin_1 => "000110010001101111", pass => false),
  (xin_0 => "001000100110001001", xin_1 => "001011111000011011", pass => false),
  (xin_0 => "001110011000001010", xin_1 => "000101100000001001", pass => false),
  (xin_0 => "001000101010111000", xin_1 => "000100111100001010", pass => true),
  (xin_0 => "001011010011000011", xin_1 => "001001000101110111", pass => false),
  (xin_0 => "001000111101101010", xin_1 => "001011111011000101", pass => false),
  (xin_0 => "000111100101010010", xin_1 => "000001100001010001", pass => false),
  (xin_0 => "000101111000100111", xin_1 => "001010110000010000", pass => false),
  (xin_0 => "001001111000011000", xin_1 => "000111000101011110", pass => true),
  (xin_0 => "001001101010101110", xin_1 => "000011011111100001", pass => false),
  (xin_0 => "001101010011110100", xin_1 => "000110000010101111", pass => false),
  (xin_0 => "001011010011100000", xin_1 => "000101110001010111", pass => true),
  (xin_0 => "001001110110101101", xin_1 => "001011100101100010", pass => false),
  (xin_0 => "001001101011001100", xin_1 => "000001110001110000", pass => false),
  (xin_0 => "001100010001001110", xin_1 => "000101111111100100", pass => false),
  (xin_0 => "001000010011101001", xin_1 => "000010010101000000", pass => false),
  (xin_0 => "001100110010100101", xin_1 => "001010010111000000", pass => true),
  (xin_0 => "000110101100111001", xin_1 => "001001111011010011", pass => false),
  (xin_0 => "000110010011000010", xin_1 => "000010111100000000", pass => false),
  (xin_0 => "000111111001011110", xin_1 => "000101111110011101", pass => true),
  (xin_0 => "000101101000100010", xin_1 => "000100100001010010", pass => true),
  (xin_0 => "000111100001000010", xin_1 => "000010111010011000", pass => false),
  (xin_0 => "000111010110010000", xin_1 => "000101000100101100", pass => true),
  (xin_0 => "000101000101100100", xin_1 => "000100010000101111", pass => true),
  (xin_0 => "000110101000000000", xin_1 => "001010000001100010", pass => false),
  (xin_0 => "001001100000100001", xin_1 => "001011011101001110", pass => false),
  (xin_0 => "000100001011111101", xin_1 => "000010010111101001", pass => true),
  (xin_0 => "001001011101100101", xin_1 => "000010110110100110", pass => false),
  (xin_0 => "001000010011011010", xin_1 => "000011001000111111", pass => false),
  (xin_0 => "001001010001000000", xin_1 => "000010100011101000", pass => false),
  (xin_0 => "001001101000100110", xin_1 => "000010111111100010", pass => false),
  (xin_0 => "001010101111110011", xin_1 => "001011001111001100", pass => false),
  (xin_0 => "001100101101011110", xin_1 => "001000100000010101", pass => false),
  (xin_0 => "001000101010011011", xin_1 => "000011000001110011", pass => false),
  (xin_0 => "001001000000010101", xin_1 => "000011001010000001", pass => false),
  (xin_0 => "001001101000111000", xin_1 => "000010011001010011", pass => false),
  (xin_0 => "000100111111100111", xin_1 => "001001000011000110", pass => false),
  (xin_0 => "000101000100111010", xin_1 => "000100111101000110", pass => true),
  (xin_0 => "001011001001111010", xin_1 => "000010101100100000", pass => true),
  (xin_0 => "000110110010011110", xin_1 => "000100101011011101", pass => true),
  (xin_0 => "001100011100011000", xin_1 => "000011110111001001", pass => true),
  (xin_0 => "000111101001111000", xin_1 => "001000111111100001", pass => false),
  (xin_0 => "001001001100001010", xin_1 => "000111011111111011", pass => true),
  (xin_0 => "001001011001100101", xin_1 => "001000001000111000", pass => true),
  (xin_0 => "001000100110000010", xin_1 => "000011010101101010", pass => false),
  (xin_0 => "000011100110001010", xin_1 => "000101001010111101", pass => true),
  (xin_0 => "001010000010110101", xin_1 => "000100010001100011", pass => true),
  (xin_0 => "001010000011000101", xin_1 => "000110000010101101", pass => true),
  (xin_0 => "000111100111100100", xin_1 => "000111010001001111", pass => true),
  (xin_0 => "000111001110000001", xin_1 => "000010000010101101", pass => false),
  (xin_0 => "001100000010001000", xin_1 => "000111000010010101", pass => false),
  (xin_0 => "001101100101111111", xin_1 => "000101101011000001", pass => false),
  (xin_0 => "010000010110010111", xin_1 => "001010011110101000", pass => true),
  (xin_0 => "001100111010100111", xin_1 => "001010101000110111", pass => true),
  (xin_0 => "001001111001011110", xin_1 => "000110001111110010", pass => true),
  (xin_0 => "000110110101010111", xin_1 => "000011011110010001", pass => false),
  (xin_0 => "001001100100000011", xin_1 => "000010010110000000", pass => false),
  (xin_0 => "001011101101101000", xin_1 => "000111100001100111", pass => false),
  (xin_0 => "001000101001011100", xin_1 => "000010110000110111", pass => false),
  (xin_0 => "000100000101011011", xin_1 => "000100100111110001", pass => true),
  (xin_0 => "001000000001010001", xin_1 => "000101001001011001", pass => true),
  (xin_0 => "001100111111001001", xin_1 => "000011100101000000", pass => true),
  (xin_0 => "001000110000001010", xin_1 => "000010010001000010", pass => false),
  (xin_0 => "001001110101101010", xin_1 => "000101101111010100", pass => true),
  (xin_0 => "001101000001000110", xin_1 => "001000110100111000", pass => false),
  (xin_0 => "001100101011100000", xin_1 => "001001011111011110", pass => false),
  (xin_0 => "001001010101110101", xin_1 => "000010101001010111", pass => false),
  (xin_0 => "000110100011110110", xin_1 => "000011010010100101", pass => false),
  (xin_0 => "000101101000010110", xin_1 => "000100010000101111", pass => true),
  (xin_0 => "000100100000010111", xin_1 => "000100110011110101", pass => true),
  (xin_0 => "001101101110111101", xin_1 => "000110010110011011", pass => false),
  (xin_0 => "000100001001000000", xin_1 => "000011110100011111", pass => true),
  (xin_0 => "000111011000001111", xin_1 => "000110001010100110", pass => true),
  (xin_0 => "000101101110010101", xin_1 => "000110001110111001", pass => true),
  (xin_0 => "001100101000110100", xin_1 => "001011000110001001", pass => true),
  (xin_0 => "000111101101001111", xin_1 => "000001111110011001", pass => false),
  (xin_0 => "001011000000101011", xin_1 => "000110011000110110", pass => true),
  (xin_0 => "001100000010100110", xin_1 => "000111011100001000", pass => false),
  (xin_0 => "000111101111000100", xin_1 => "001001100110110111", pass => false),
  (xin_0 => "001100101100100110", xin_1 => "001000000111100001", pass => false),
  (xin_0 => "001010101010010011", xin_1 => "001000011001100011", pass => false),
  (xin_0 => "000111010100001001", xin_1 => "000101111110100100", pass => true),
  (xin_0 => "001010010000010100", xin_1 => "001000001100100101", pass => false),
  (xin_0 => "001010000010010001", xin_1 => "001010101110000101", pass => false),
  (xin_0 => "001011111000010111", xin_1 => "000011010111101010", pass => true),
  (xin_0 => "001010001010011101", xin_1 => "000100000100010001", pass => true),
  (xin_0 => "001000010001111001", xin_1 => "000101000111110010", pass => true),
  (xin_0 => "000011101110011000", xin_1 => "000111110101011111", pass => false),
  (xin_0 => "010000010001011110", xin_1 => "001010110001111101", pass => true),
  (xin_0 => "001010110100010010", xin_1 => "000101001010010110", pass => true),
  (xin_0 => "000111100011010001", xin_1 => "000010100101010010", pass => false),
  (xin_0 => "001011101011011101", xin_1 => "001001110000001111", pass => false),
  (xin_0 => "000101001101100101", xin_1 => "000010110001001110", pass => true),
  (xin_0 => "001011111010000111", xin_1 => "001001010000100000", pass => false),
  (xin_0 => "001000100011101011", xin_1 => "001010100101111010", pass => false),
  (xin_0 => "001000111000000111", xin_1 => "000011010101011011", pass => false),
  (xin_0 => "001001101111101001", xin_1 => "000001110100110110", pass => false),
  (xin_0 => "001100110000101011", xin_1 => "000110100101011110", pass => false),
  (xin_0 => "000111000010111101", xin_1 => "000111111010011100", pass => true),
  (xin_0 => "000100101001001111", xin_1 => "000101100011100101", pass => true),
  (xin_0 => "001001010100010000", xin_1 => "001100110010101111", pass => false),
  (xin_0 => "000111111011000011", xin_1 => "000010101100111100", pass => false),
  (xin_0 => "001001110010101111", xin_1 => "000100101010011100", pass => true),
  (xin_0 => "001011101001111111", xin_1 => "000010011110000111", pass => true),
  (xin_0 => "000110011111001111", xin_1 => "000010011000111111", pass => false),
  (xin_0 => "001000111001000111", xin_1 => "000010111011001111", pass => false),
  (xin_0 => "000011111111111100", xin_1 => "000010010010101010", pass => true),
  (xin_0 => "000101001101101111", xin_1 => "001010110111001010", pass => false),
  (xin_0 => "000111011111000100", xin_1 => "001001111111111010", pass => false),
  (xin_0 => "001001101111010101", xin_1 => "000100011011100011", pass => true),
  (xin_0 => "001010101110010000", xin_1 => "001000001100110111", pass => false),
  (xin_0 => "001100100110110110", xin_1 => "000111101000011011", pass => false),
  (xin_0 => "001011100100001101", xin_1 => "001001000110101101", pass => false),
  (xin_0 => "001110110111001011", xin_1 => "001010010111110000", pass => true),
  (xin_0 => "000100010111011001", xin_1 => "000011101010110101", pass => true),
  (xin_0 => "000100110010011111", xin_1 => "000100101100010111", pass => true),
  (xin_0 => "000110100100101100", xin_1 => "000001110101110100", pass => false),
  (xin_0 => "001010010100100000", xin_1 => "001010011001001100", pass => false),
  (xin_0 => "000110100101110101", xin_1 => "001001110011010111", pass => false),
  (xin_0 => "001011100000001111", xin_1 => "000111000100000000", pass => false),
  (xin_0 => "001000101010000101", xin_1 => "000101110101001111", pass => true),
  (xin_0 => "001100010110100000", xin_1 => "000010000000010101", pass => true),
  (xin_0 => "000100111001111000", xin_1 => "000111111010000111", pass => false),
  (xin_0 => "000110000110001110", xin_1 => "000010010110111010", pass => false),
  (xin_0 => "001000000000100000", xin_1 => "000110101111010101", pass => true),
  (xin_0 => "000101110110010010", xin_1 => "000100010101101000", pass => true),
  (xin_0 => "001010001000011101", xin_1 => "000011010111110000", pass => false),
  (xin_0 => "000111001100011001", xin_1 => "000011100000100100", pass => false),
  (xin_0 => "001010010011111110", xin_1 => "001100000001111001", pass => false),
  (xin_0 => "001100000001100011", xin_1 => "001000100011000100", pass => false),
  (xin_0 => "001000111110100101", xin_1 => "001010001101010100", pass => false),
  (xin_0 => "001001010001010101", xin_1 => "000111111010001111", pass => true),
  (xin_0 => "001110001100000100", xin_1 => "000100100011011011", pass => false),
  (xin_0 => "001101111101100100", xin_1 => "001010000011111011", pass => true),
  (xin_0 => "001000100110100100", xin_1 => "000011000010100010", pass => false),
  (xin_0 => "001011011000110110", xin_1 => "001010100011011101", pass => false),
  (xin_0 => "001110000001000110", xin_1 => "000110010001101011", pass => false),
  (xin_0 => "001001100011011100", xin_1 => "000010000001111000", pass => false),
  (xin_0 => "001011001101110100", xin_1 => "001000111111110100", pass => false),
  (xin_0 => "001100110010101111", xin_1 => "001011001011000001", pass => true),
  (xin_0 => "001000000010110001", xin_1 => "000100000010100011", pass => false),
  (xin_0 => "000101001001001100", xin_1 => "000110110000101100", pass => true),
  (xin_0 => "001011000111010110", xin_1 => "001001001111010100", pass => false),
  (xin_0 => "000111010100110010", xin_1 => "000011100100101011", pass => false),
  (xin_0 => "000110100000010100", xin_1 => "000101000101001001", pass => true),
  (xin_0 => "001000110000000110", xin_1 => "000011100000001111", pass => false),
  (xin_0 => "000111100001010011", xin_1 => "000100000010100111", pass => false),
  (xin_0 => "001001110100011010", xin_1 => "001010111101111110", pass => false),
  (xin_0 => "000110111101011011", xin_1 => "000010110001001010", pass => false),
  (xin_0 => "001100111100000100", xin_1 => "000000111011011011", pass => true),
  (xin_0 => "001001111000110001", xin_1 => "000011000100110001", pass => false),
  (xin_0 => "001000010110101101", xin_1 => "000100110010010110", pass => true),
  (xin_0 => "001010111001000100", xin_1 => "001001001101010011", pass => false),
  (xin_0 => "001110010100111010", xin_1 => "001011000110111100", pass => true),
  (xin_0 => "001001010111101010", xin_1 => "001010111110011001", pass => false),
  (xin_0 => "001000001110000110", xin_1 => "000100111111100011", pass => true),
  (xin_0 => "001101000001101001", xin_1 => "001000000100100110", pass => false),
  (xin_0 => "001010000101100100", xin_1 => "000101111101000010", pass => true),
  (xin_0 => "000111110111001111", xin_1 => "001010010001110110", pass => false),
  (xin_0 => "000111000110100001", xin_1 => "001010000111110010", pass => false),
  (xin_0 => "001000101001010100", xin_1 => "000011011001000011", pass => false),
  (xin_0 => "000111010000001001", xin_1 => "001001010011001001", pass => false),
  (xin_0 => "000111100001111011", xin_1 => "000100111011000100", pass => true),
  (xin_0 => "001001001001110110", xin_1 => "000011101101100100", pass => false),
  (xin_0 => "001100010100000001", xin_1 => "001000100101100101", pass => false),
  (xin_0 => "000111101001001100", xin_1 => "000010100001000110", pass => false),
  (xin_0 => "001011001110110101", xin_1 => "001010001100100011", pass => false),
  (xin_0 => "001001001001111101", xin_1 => "000010011010100000", pass => false),
  (xin_0 => "001010001000110010", xin_1 => "000110110111110010", pass => true),
  (xin_0 => "001001101101110001", xin_1 => "000001101111000100", pass => false),
  (xin_0 => "001000001110100010", xin_1 => "001000110011000111", pass => true),
  (xin_0 => "001100001000110001", xin_1 => "001000000100000010", pass => false),
  (xin_0 => "001000101000000011", xin_1 => "001000001000010100", pass => true),
  (xin_0 => "001010000001100000", xin_1 => "001011011000000000", pass => false),
  (xin_0 => "000111000111010111", xin_1 => "000010101111101110", pass => false),
  (xin_0 => "001001110101111010", xin_1 => "000110100101111110", pass => true),
  (xin_0 => "000011111010010010", xin_1 => "001000010101010101", pass => false),
  (xin_0 => "001000010111011110", xin_1 => "001011001101100000", pass => false),
  (xin_0 => "001100011010010111", xin_1 => "000111111010011000", pass => false),
  (xin_0 => "001000111100100001", xin_1 => "000011001000100010", pass => false),
  (xin_0 => "001100100110100101", xin_1 => "000011000110111101", pass => true),
  (xin_0 => "000111111101110110", xin_1 => "001010111011101001", pass => false),
  (xin_0 => "000100110100101101", xin_1 => "000101001001001100", pass => true),
  (xin_0 => "000100110111111101", xin_1 => "001001100010001110", pass => false),
  (xin_0 => "000100010101010110", xin_1 => "001001000000001110", pass => false),
  (xin_0 => "000011000100101110", xin_1 => "000111010100011011", pass => false),
  (xin_0 => "001100100100011110", xin_1 => "000101100111001011", pass => false),
  (xin_0 => "001101011000110111", xin_1 => "000011000001110101", pass => true),
  (xin_0 => "000101111000000101", xin_1 => "000100100011110100", pass => true),
  (xin_0 => "000100010110101011", xin_1 => "000011111001100111", pass => true),
  (xin_0 => "001010010000010000", xin_1 => "000110000101000011", pass => true),
  (xin_0 => "000111100010101001", xin_1 => "000100100110010110", pass => true),
  (xin_0 => "000011100110111011", xin_1 => "000110100000101100", pass => false),
  (xin_0 => "000111101110111100", xin_1 => "000010111010101111", pass => false),
  (xin_0 => "000110100010100100", xin_1 => "000010011111001011", pass => false),
  (xin_0 => "000110110001010001", xin_1 => "001001100101100001", pass => false),
  (xin_0 => "001000110000000011", xin_1 => "000010100100101101", pass => false),
  (xin_0 => "001000001100101001", xin_1 => "000110110110010001", pass => true),
  (xin_0 => "000110101011000110", xin_1 => "000101111000100010", pass => true),
  (xin_0 => "001100110111101101", xin_1 => "001000001011111001", pass => false),
  (xin_0 => "001011010100010011", xin_1 => "000101110100101100", pass => true),
  (xin_0 => "001100001000100101", xin_1 => "001000000100000101", pass => false),
  (xin_0 => "001000101111001111", xin_1 => "000010000001111001", pass => false),
  (xin_0 => "001100011100011011", xin_1 => "000101100101001010", pass => false),
  (xin_0 => "001101011111100110", xin_1 => "000111101100100111", pass => false),
  (xin_0 => "000101100100001010", xin_1 => "001001100000111011", pass => false),
  (xin_0 => "001001000100010100", xin_1 => "000010000111101101", pass => false),
  (xin_0 => "000111110010111111", xin_1 => "001010001100001011", pass => false),
  (xin_0 => "000110111110000000", xin_1 => "000111100111111100", pass => true),
  (xin_0 => "000111001001001011", xin_1 => "001011001111011001", pass => false),
  (xin_0 => "000110100110000001", xin_1 => "000110111011010010", pass => true),
  (xin_0 => "001000000100011111", xin_1 => "000110111110101000", pass => true),
  (xin_0 => "001011111111100001", xin_1 => "000111100100111101", pass => false),
  (xin_0 => "000111001110010101", xin_1 => "000110111011110001", pass => true),
  (xin_0 => "001000100110010100", xin_1 => "000011110001010111", pass => false),
  (xin_0 => "001011001101110111", xin_1 => "000111011111010111", pass => false),
  (xin_0 => "000011011111011011", xin_1 => "000100000001001110", pass => true),
  (xin_0 => "001000111111000111", xin_1 => "000001110011010001", pass => false),
  (xin_0 => "001001011000101010", xin_1 => "000101010101001100", pass => true),
  (xin_0 => "000111100101011001", xin_1 => "000111011110100110", pass => true),
  (xin_0 => "000110010000100010", xin_1 => "001000100010000010", pass => false),
  (xin_0 => "001011010101011111", xin_1 => "000110110011111001", pass => false),
  (xin_0 => "001001010000001000", xin_1 => "000111001110101010", pass => true),
  (xin_0 => "000111010010011111", xin_1 => "001010001110011101", pass => false),
  (xin_0 => "001001000011001110", xin_1 => "000111001101010110", pass => true),
  (xin_0 => "001011000101111110", xin_1 => "000110101001101010", pass => true),
  (xin_0 => "001000100111100000", xin_1 => "001010000100000000", pass => false),
  (xin_0 => "000111001001000000", xin_1 => "001010011010010001", pass => false),
  (xin_0 => "001010011001100111", xin_1 => "000010101010100100", pass => false),
  (xin_0 => "001011011111100000", xin_1 => "000011010010000010", pass => true),
  (xin_0 => "000101110101111110", xin_1 => "001001110001000001", pass => false),
  (xin_0 => "000011110011000001", xin_1 => "000100011101010101", pass => true),
  (xin_0 => "000100100100000010", xin_1 => "000011001101011100", pass => true),
  (xin_0 => "001000100111011011", xin_1 => "000010000110001000", pass => false),
  (xin_0 => "000111011100110100", xin_1 => "000011110011001101", pass => false),
  (xin_0 => "000011100111101011", xin_1 => "000011100110001110", pass => true),
  (xin_0 => "000101001001010101", xin_1 => "000101100010000000", pass => true),
  (xin_0 => "001100101010000010", xin_1 => "000111010111001101", pass => false),
  (xin_0 => "001011100100110001", xin_1 => "000011001101001011", pass => true),
  (xin_0 => "001001001101111101", xin_1 => "000111101110100100", pass => true),
  (xin_0 => "000110110001011001", xin_1 => "001001100100010100", pass => false),
  (xin_0 => "000110100011010010", xin_1 => "001001011101010110", pass => false),
  (xin_0 => "001110010101011100", xin_1 => "000101100101001101", pass => false),
  (xin_0 => "000100011101010101", xin_1 => "000100001101100111", pass => true),
  (xin_0 => "001001110110001100", xin_1 => "000011000001001010", pass => false),
  (xin_0 => "001011000000001001", xin_1 => "000011110111001111", pass => true),
  (xin_0 => "001001111110100100", xin_1 => "000010100111010111", pass => false),
  (xin_0 => "001011000011101001", xin_1 => "000111000110101101", pass => false),
  (xin_0 => "000110111111110101", xin_1 => "001001110100010011", pass => false),
  (xin_0 => "001100101011101001", xin_1 => "000010100111000111", pass => true),
  (xin_0 => "000101011001110111", xin_1 => "001000110000001100", pass => false),
  (xin_0 => "001001100010110001", xin_1 => "000011000000101101", pass => false),
  (xin_0 => "000101000111000001", xin_1 => "001001011111111101", pass => false),
  (xin_0 => "001011101101100001", xin_1 => "000011110110011010", pass => true),
  (xin_0 => "000110101011010111", xin_1 => "000101001000010001", pass => true),
  (xin_0 => "010000100011001000", xin_1 => "001001100111101011", pass => true),
  (xin_0 => "001001001110010101", xin_1 => "001100100110110011", pass => false),
  (xin_0 => "000101000001111111", xin_1 => "000100011111101010", pass => true),
  (xin_0 => "001011111001100001", xin_1 => "000110011001000101", pass => false),
  (xin_0 => "001011111010111101", xin_1 => "000101001010010000", pass => true),
  (xin_0 => "001000010111101111", xin_1 => "001010010101000000", pass => false),
  (xin_0 => "001001011011101101", xin_1 => "000010011011101000", pass => false),
  (xin_0 => "000111111100000011", xin_1 => "001100100000010111", pass => false),
  (xin_0 => "001011111000110001", xin_1 => "000101100110101110", pass => true),
  (xin_0 => "000110100010010001", xin_1 => "001010101111001110", pass => false),
  (xin_0 => "000100000010000100", xin_1 => "000000110010010001", pass => true),
  (xin_0 => "000100100110011010", xin_1 => "000110011111000010", pass => true),
  (xin_0 => "000110010111111111", xin_1 => "000010101011010000", pass => false),
  (xin_0 => "001100011110110101", xin_1 => "000111100000111100", pass => false),
  (xin_0 => "001000101100110000", xin_1 => "000111000000001010", pass => true),
  (xin_0 => "000011110010001111", xin_1 => "000100011000011001", pass => true),
  (xin_0 => "001001101110001100", xin_1 => "001010011111011101", pass => false),
  (xin_0 => "001010101001100101", xin_1 => "001001101110010110", pass => false),
  (xin_0 => "000111101001111000", xin_1 => "000101001001101011", pass => true),
  (xin_0 => "000111011011010000", xin_1 => "001000111011000100", pass => false),
  (xin_0 => "000100011101010110", xin_1 => "001000010101101101", pass => false),
  (xin_0 => "001000101011001010", xin_1 => "000110110011011101", pass => true),
  (xin_0 => "001000010101001000", xin_1 => "000011001010110111", pass => false),
  (xin_0 => "001100100101111110", xin_1 => "000011011101001100", pass => true),
  (xin_0 => "001000110111001100", xin_1 => "000011001001010010", pass => false),
  (xin_0 => "000111001001010100", xin_1 => "001011100011010100", pass => false),
  (xin_0 => "000101111100100100", xin_1 => "001001001101111101", pass => false),
  (xin_0 => "000110011010001001", xin_1 => "000010101100101000", pass => false),
  (xin_0 => "001100100110101110", xin_1 => "000110101010101011", pass => false),
  (xin_0 => "000111110011100110", xin_1 => "000010000001111011", pass => false),
  (xin_0 => "001011001000100111", xin_1 => "001011110011111001", pass => false),
  (xin_0 => "001000001010001100", xin_1 => "000111101101101110", pass => true),
  (xin_0 => "001001000100100111", xin_1 => "000010110010011111", pass => false),
  (xin_0 => "000101110111111100", xin_1 => "000110110001110010", pass => true),
  (xin_0 => "001001011010000101", xin_1 => "000011011000110101", pass => false),
  (xin_0 => "000011000000110011", xin_1 => "000000010111110000", pass => true),
  (xin_0 => "000111111100011101", xin_1 => "000110100101100111", pass => true),
  (xin_0 => "000011001000000110", xin_1 => "000111100011111110", pass => false),
  (xin_0 => "001000000101000100", xin_1 => "000101111000000100", pass => true),
  (xin_0 => "000111000011100010", xin_1 => "000001110110011101", pass => false),
  (xin_0 => "000011000111110010", xin_1 => "000000100111100101", pass => true),
  (xin_0 => "001011110011001011", xin_1 => "000100110110101110", pass => true),
  (xin_0 => "000110101100110111", xin_1 => "000010001011101010", pass => false),
  (xin_0 => "001100110101011101", xin_1 => "001010011000001101", pass => true),
  (xin_0 => "001001010011011011", xin_1 => "000110111001000111", pass => true),
  (xin_0 => "000101101000111100", xin_1 => "001000110011101010", pass => false),
  (xin_0 => "000101110101011011", xin_1 => "001000011010101110", pass => false),
  (xin_0 => "001000100001010101", xin_1 => "000010100100111000", pass => false),
  (xin_0 => "001000100010110000", xin_1 => "000110111011100100", pass => true),
  (xin_0 => "000111111110100001", xin_1 => "001011110111000111", pass => false),
  (xin_0 => "000111100100111110", xin_1 => "000011001000011011", pass => false),
  (xin_0 => "001000011110111001", xin_1 => "000101001101100011", pass => true),
  (xin_0 => "000111101011111001", xin_1 => "000011001111001000", pass => false),
  (xin_0 => "000111110111000111", xin_1 => "000011010001010101", pass => false),
  (xin_0 => "001000101110011100", xin_1 => "000010101101000001", pass => false),
  (xin_0 => "000101111111011111", xin_1 => "000010101000111110", pass => false),
  (xin_0 => "001100101101101010", xin_1 => "000110110010110011", pass => false),
  (xin_0 => "001011001110101010", xin_1 => "000110010111111011", pass => true),
  (xin_0 => "001000111010101000", xin_1 => "000010010111101000", pass => false),
  (xin_0 => "001100100000100001", xin_1 => "000101111000010001", pass => false),
  (xin_0 => "001000100001111101", xin_1 => "000110101000010010", pass => true),
  (xin_0 => "001001101011101111", xin_1 => "000101000010111000", pass => true),
  (xin_0 => "001111101011001010", xin_1 => "001010001010110000", pass => true),
  (xin_0 => "000111000110010101", xin_1 => "001000010111110100", pass => true),
  (xin_0 => "001000000000000101", xin_1 => "000011100111101000", pass => false),
  (xin_0 => "000110001000011010", xin_1 => "000111110001111111", pass => true),
  (xin_0 => "001110000000011000", xin_1 => "000111111110110000", pass => false),
  (xin_0 => "001101001001110011", xin_1 => "000010011011000010", pass => true),
  (xin_0 => "001011101110011011", xin_1 => "000110100001101111", pass => false),
  (xin_0 => "001011110010000011", xin_1 => "000010000000110010", pass => true),
  (xin_0 => "001010000000111001", xin_1 => "000110101110100001", pass => true),
  (xin_0 => "000011011111011111", xin_1 => "000011010000000100", pass => true),
  (xin_0 => "001011110100100101", xin_1 => "001000100100100000", pass => false),
  (xin_0 => "000110001001110001", xin_1 => "001001111100110001", pass => false),
  (xin_0 => "001000100011010011", xin_1 => "000101000111111110", pass => true),
  (xin_0 => "000101001011000110", xin_1 => "000011101101001111", pass => true),
  (xin_0 => "000111010101000110", xin_1 => "000010110100011011", pass => false),
  (xin_0 => "001101111110101000", xin_1 => "001001001101000101", pass => true),
  (xin_0 => "001001011111011000", xin_1 => "000111000001010010", pass => true),
  (xin_0 => "001011100011111011", xin_1 => "000010000101000111", pass => true),
  (xin_0 => "000101010110001010", xin_1 => "000110001100100010", pass => true),
  (xin_0 => "001011110001100101", xin_1 => "001000111001010001", pass => false),
  (xin_0 => "000111011101110011", xin_1 => "001010001001001001", pass => false),
  (xin_0 => "000110111011110000", xin_1 => "001010010100011000", pass => false),
  (xin_0 => "001000010111010100", xin_1 => "000010111101000001", pass => false),
  (xin_0 => "000110010110001000", xin_1 => "001010110000011111", pass => false),
  (xin_0 => "001010001111000101", xin_1 => "001010111010110011", pass => false),
  (xin_0 => "001001111011001011", xin_1 => "001100010001110001", pass => false),
  (xin_0 => "000101001111100110", xin_1 => "001000011010101010", pass => false),
  (xin_0 => "000100110011111111", xin_1 => "001000011000000111", pass => false),
  (xin_0 => "000111101101000111", xin_1 => "001001111001000010", pass => false),
  (xin_0 => "001100000001110100", xin_1 => "000100110110100010", pass => true),
  (xin_0 => "001101110000110101", xin_1 => "001000010001010011", pass => false),
  (xin_0 => "001011101011110010", xin_1 => "000110111110110001", pass => false),
  (xin_0 => "001111010110110100", xin_1 => "001001111001011001", pass => true),
  (xin_0 => "000110100011000000", xin_1 => "001001001111101001", pass => false),
  (xin_0 => "000110100001100001", xin_1 => "000111010011110111", pass => true),
  (xin_0 => "000011101010001100", xin_1 => "000111011000001101", pass => false),
  (xin_0 => "000011101011001100", xin_1 => "001000111110010111", pass => false),
  (xin_0 => "001101010011010011", xin_1 => "000110010111001010", pass => false),
  (xin_0 => "001011000000001000", xin_1 => "001010011001100011", pass => false),
  (xin_0 => "000111111000100000", xin_1 => "000011010010110101", pass => false),
  (xin_0 => "000111011010111000", xin_1 => "000111010101101001", pass => true),
  (xin_0 => "001000010100110111", xin_1 => "000010000001110010", pass => false),
  (xin_0 => "000101110000011010", xin_1 => "000010110010111101", pass => false),
  (xin_0 => "001101000111100010", xin_1 => "000000111110011011", pass => true),
  (xin_0 => "001110001000111000", xin_1 => "000100110101010100", pass => false),
  (xin_0 => "000110001011011101", xin_1 => "000110010110001010", pass => true),
  (xin_0 => "001011101001100011", xin_1 => "000101000101100111", pass => true),
  (xin_0 => "000110011010000110", xin_1 => "000001110010110110", pass => false),
  (xin_0 => "000110010111100010", xin_1 => "001010000001011111", pass => false),
  (xin_0 => "000110100001111110", xin_1 => "000010000110101001", pass => false),
  (xin_0 => "001000111100011001", xin_1 => "000101111111011101", pass => true),
  (xin_0 => "001000000110111101", xin_1 => "000011100111100100", pass => false),
  (xin_0 => "000100011110111110", xin_1 => "000100010001011001", pass => true),
  (xin_0 => "001000000101101100", xin_1 => "000010101100100000", pass => false),
  (xin_0 => "001010001111011111", xin_1 => "000110101000110101", pass => true),
  (xin_0 => "000111010111101100", xin_1 => "000111100100100111", pass => true),
  (xin_0 => "001000011001110110", xin_1 => "000110101111001110", pass => true),
  (xin_0 => "001000001000000100", xin_1 => "000010111000011010", pass => false),
  (xin_0 => "001001101010100111", xin_1 => "000011111001011001", pass => false),
  (xin_0 => "000110101000000111", xin_1 => "000010111010110101", pass => false),
  (xin_0 => "000100100001010000", xin_1 => "000111101111111100", pass => false),
  (xin_0 => "000101111011110101", xin_1 => "000001111010100100", pass => false),
  (xin_0 => "001001110010111011", xin_1 => "001010010010111101", pass => false),
  (xin_0 => "001001001010110100", xin_1 => "001001011000010111", pass => false),
  (xin_0 => "001010100000101100", xin_1 => "000010000000111001", pass => false),
  (xin_0 => "000101001010011010", xin_1 => "000101010000001111", pass => true),
  (xin_0 => "000001100001110011", xin_1 => "000101111111010100", pass => false),
  (xin_0 => "000111001101111100", xin_1 => "000100101001001011", pass => true),
  (xin_0 => "000010100110110010", xin_1 => "000010010001100101", pass => true),
  (xin_0 => "000100010111110100", xin_1 => "000111100111010000", pass => false),
  (xin_0 => "000011100010001010", xin_1 => "000100100010100000", pass => true),
  (xin_0 => "000101001001110010", xin_1 => "000100010100100110", pass => true),
  (xin_0 => "001100010100110101", xin_1 => "000010011100110100", pass => true),
  (xin_0 => "000110110111110110", xin_1 => "000010011010100100", pass => false),
  (xin_0 => "000100011000110111", xin_1 => "000010011010000010", pass => true),
  (xin_0 => "000110011010000001", xin_1 => "000111101111101011", pass => true),
  (xin_0 => "001101011011010110", xin_1 => "001011100011011100", pass => true),
  (xin_0 => "000101101101011100", xin_1 => "000101010001010011", pass => true),
  (xin_0 => "001100100011111111", xin_1 => "000111111010100111", pass => false),
  (xin_0 => "001000010100011000", xin_1 => "000111110100011101", pass => true),
  (xin_0 => "001101001000010111", xin_1 => "001000111101010100", pass => false),
  (xin_0 => "001010000111111001", xin_1 => "000110010000100000", pass => true),
  (xin_0 => "001100010000010111", xin_1 => "000111010111101111", pass => false),
  (xin_0 => "001110000000000100", xin_1 => "000110110100011100", pass => false),
  (xin_0 => "001001101111101011", xin_1 => "001011010100011110", pass => false),
  (xin_0 => "000110001101000101", xin_1 => "001001010001101000", pass => false),
  (xin_0 => "001001001010101000", xin_1 => "000011001010000100", pass => false),
  (xin_0 => "000100000101110110", xin_1 => "000100101011011001", pass => true),
  (xin_0 => "001011110001101101", xin_1 => "000010001100110100", pass => true),
  (xin_0 => "000111001001111001", xin_1 => "001010110111001000", pass => false),
  (xin_0 => "000010111110101000", xin_1 => "000010011111010000", pass => true),
  (xin_0 => "000011010101100001", xin_1 => "000011000101111110", pass => true),
  (xin_0 => "001011100111010000", xin_1 => "001000101110001000", pass => false),
  (xin_0 => "001011011010110001", xin_1 => "001000000010110100", pass => false),
  (xin_0 => "001000101000000111", xin_1 => "000101101000001110", pass => true),
  (xin_0 => "001001100111101001", xin_1 => "000010101110101100", pass => false),
  (xin_0 => "001001000010000100", xin_1 => "000100001001101100", pass => false),
  (xin_0 => "001001011101101100", xin_1 => "001100000111101101", pass => false),
  (xin_0 => "000111000001100011", xin_1 => "000010001001100100", pass => false),
  (xin_0 => "000111010011101101", xin_1 => "000011100100110100", pass => false),
  (xin_0 => "000011100111100010", xin_1 => "000011010100001010", pass => true),
  (xin_0 => "001001101111000010", xin_1 => "000110011000000111", pass => true),
  (xin_0 => "000111011000100111", xin_1 => "000101001110000001", pass => true),
  (xin_0 => "001110110110000001", xin_1 => "001001100101011110", pass => true),
  (xin_0 => "001010010100000111", xin_1 => "000011111001110100", pass => true),
  (xin_0 => "000101110110111111", xin_1 => "001001001001110110", pass => false),
  (xin_0 => "001000101001111011", xin_1 => "000001000001000110", pass => false),
  (xin_0 => "001001110010100000", xin_1 => "001011001001111010", pass => false),
  (xin_0 => "000111101000101010", xin_1 => "000010010010000111", pass => false),
  (xin_0 => "001010110111001001", xin_1 => "001001000000001100", pass => false),
  (xin_0 => "001100110110000101", xin_1 => "000111001100111010", pass => false),
  (xin_0 => "001000010100100101", xin_1 => "001100100101001010", pass => false),
  (xin_0 => "001101001001000110", xin_1 => "000111000011100110", pass => false),
  (xin_0 => "000100001000000011", xin_1 => "000011100100010000", pass => true),
  (xin_0 => "000111110010000010", xin_1 => "000110110001001111", pass => true),
  (xin_0 => "001100000011010101", xin_1 => "000010000001101110", pass => true),
  (xin_0 => "001000101110110100", xin_1 => "000010110100111100", pass => false),
  (xin_0 => "001010110100101111", xin_1 => "001001111110011101", pass => false),
  (xin_0 => "001000100010000011", xin_1 => "001011010100001010", pass => false),
  (xin_0 => "001010010011111100", xin_1 => "000101010000001010", pass => true),
  (xin_0 => "001011001110000001", xin_1 => "001011101100001100", pass => false),
  (xin_0 => "001000111101010100", xin_1 => "000111000001100110", pass => true),
  (xin_0 => "000100000111101101", xin_1 => "001001100101000100", pass => false),
  (xin_0 => "001001011100100011", xin_1 => "000100000010100111", pass => false),
  (xin_0 => "001011110001100011", xin_1 => "000011010101100100", pass => true),
  (xin_0 => "001010100110110010", xin_1 => "001010100010000000", pass => false),
  (xin_0 => "001100000101011001", xin_1 => "001001010111101101", pass => false),
  (xin_0 => "000110011001011011", xin_1 => "000100011101010110", pass => true),
  (xin_0 => "001000100011010100", xin_1 => "000010011000010100", pass => false),
  (xin_0 => "000110010110010010", xin_1 => "000010011011111010", pass => false),
  (xin_0 => "001011010111000100", xin_1 => "001010010100101100", pass => false),
  (xin_0 => "001101001111000110", xin_1 => "000011000001111101", pass => true),
  (xin_0 => "001011011001000101", xin_1 => "000001111101001000", pass => true),
  (xin_0 => "000010110001101000", xin_1 => "000101001011001000", pass => true),
  (xin_0 => "000101001000000010", xin_1 => "000101000000001110", pass => true),
  (xin_0 => "000111101011011110", xin_1 => "001001111100110000", pass => false),
  (xin_0 => "000110000000101010", xin_1 => "000110001000100100", pass => true),
  (xin_0 => "000110111111001100", xin_1 => "001011000110010011", pass => false),
  (xin_0 => "001001111101111101", xin_1 => "001000111011100000", pass => false),
  (xin_0 => "001111010100100110", xin_1 => "001001000100100011", pass => true),
  (xin_0 => "001000001101111010", xin_1 => "000010010111111000", pass => false),
  (xin_0 => "000100101111100101", xin_1 => "000010011011001111", pass => true),
  (xin_0 => "001000010111001000", xin_1 => "000101101011010011", pass => true),
  (xin_0 => "001010111111000000", xin_1 => "000110010011001011", pass => true),
  (xin_0 => "001010100001111011", xin_1 => "001010100000111110", pass => false),
  (xin_0 => "000110010000100100", xin_1 => "000011100000011101", pass => false),
  (xin_0 => "001010001010100111", xin_1 => "000011100000000111", pass => true),
  (xin_0 => "001100001000000101", xin_1 => "000111100111101000", pass => false),
  (xin_0 => "000111001010101000", xin_1 => "000011110100100100", pass => false),
  (xin_0 => "000111110000110111", xin_1 => "000001111100110010", pass => false),
  (xin_0 => "000111011110101010", xin_1 => "000001111100101110", pass => false),
  (xin_0 => "001000101001000111", xin_1 => "000001101010111100", pass => false),
  (xin_0 => "001011101111011010", xin_1 => "001000110100000011", pass => false),
  (xin_0 => "000110000101000101", xin_1 => "001010011101111110", pass => false),
  (xin_0 => "001001011101011100", xin_1 => "000011100001111101", pass => false),
  (xin_0 => "000111011110110101", xin_1 => "000001000011111111", pass => false),
  (xin_0 => "001011101100111110", xin_1 => "000111100000101111", pass => false),
  (xin_0 => "000110110111010101", xin_1 => "001001110101011100", pass => false),
  (xin_0 => "001011000001010100", xin_1 => "001001010100110001", pass => false),
  (xin_0 => "000111101010011010", xin_1 => "000010011101111111", pass => false),
  (xin_0 => "001000101010110010", xin_1 => "000111011011010110", pass => true),
  (xin_0 => "000110001011001110", xin_1 => "001001011110111001", pass => false),
  (xin_0 => "000101000010011100", xin_1 => "001010001111000111", pass => false),
  (xin_0 => "001100010111101110", xin_1 => "001001000000001000", pass => false),
  (xin_0 => "001011101111010001", xin_1 => "000010001011110000", pass => true),
  (xin_0 => "001100110000111111", xin_1 => "000010011110101010", pass => true),
  (xin_0 => "000100100001100101", xin_1 => "001000101001010011", pass => false),
  (xin_0 => "000111011010110010", xin_1 => "000110100010001001", pass => true),
  (xin_0 => "001100101100101101", xin_1 => "000110111011011001", pass => false),
  (xin_0 => "001010010010111101", xin_1 => "000010010110011110", pass => false),
  (xin_0 => "001011101110011010", xin_1 => "000011110101100111", pass => true),
  (xin_0 => "001011011101100101", xin_1 => "001000000101101010", pass => false),
  (xin_0 => "001000001101110100", xin_1 => "000111011101000000", pass => true),
  (xin_0 => "001001101111111100", xin_1 => "000011001110100000", pass => false),
  (xin_0 => "001010011010100110", xin_1 => "001010101000000111", pass => false),
  (xin_0 => "000110001000110101", xin_1 => "000010111111101001", pass => false),
  (xin_0 => "001000100110101011", xin_1 => "000010100010000100", pass => false),
  (xin_0 => "001110010101100111", xin_1 => "000101001000100000", pass => false),
  (xin_0 => "001011010111111100", xin_1 => "001010000000110001", pass => false),
  (xin_0 => "000110011100101011", xin_1 => "000010110111110001", pass => false),
  (xin_0 => "001010110111001000", xin_1 => "000110000011011111", pass => true),
  (xin_0 => "000111110100010001", xin_1 => "000010011000010011", pass => false),
  (xin_0 => "000101010010101110", xin_1 => "000101010100111111", pass => true),
  (xin_0 => "001011010110010000", xin_1 => "001000110001111100", pass => false),
  (xin_0 => "000110101110110110", xin_1 => "000010100101010000", pass => false),
  (xin_0 => "000100010000111111", xin_1 => "000100000100001000", pass => true),
  (xin_0 => "001101001011000101", xin_1 => "001000001101010010", pass => false),
  (xin_0 => "001000100000000010", xin_1 => "000010101100001100", pass => false),
  (xin_0 => "000100001101000111", xin_1 => "000111111101111011", pass => false),
  (xin_0 => "000011101101000111", xin_1 => "000010100010111100", pass => true),
  (xin_0 => "001001000100011111", xin_1 => "000001101001101010", pass => false),
  (xin_0 => "000101011110101111", xin_1 => "000001111110001001", pass => false),
  (xin_0 => "001010000001000011", xin_1 => "000100110110110011", pass => true),
  (xin_0 => "001010000100101000", xin_1 => "001010111011111110", pass => false),
  (xin_0 => "001011010011001011", xin_1 => "001100000110010000", pass => false),
  (xin_0 => "001001000110111001", xin_1 => "000011001000011100", pass => false),
  (xin_0 => "001000011001010011", xin_1 => "001001011000100111", pass => false),
  (xin_0 => "001101011111011001", xin_1 => "000101000010111010", pass => false),
  (xin_0 => "001010101110110011", xin_1 => "000101101111111110", pass => true),
  (xin_0 => "001000100010000110", xin_1 => "000111101010010010", pass => true),
  (xin_0 => "001100001111011000", xin_1 => "000000111011000011", pass => true),
  (xin_0 => "001000110111111001", xin_1 => "000100011101010100", pass => true),
  (xin_0 => "000101101111011001", xin_1 => "000100111001000001", pass => true),
  (xin_0 => "000111101101100010", xin_1 => "001001101001101010", pass => false),
  (xin_0 => "000110011010000100", xin_1 => "000011010000110011", pass => false),
  (xin_0 => "001001010110010011", xin_1 => "000010000101010011", pass => false),
  (xin_0 => "001100010011111000", xin_1 => "001001011011000101", pass => false),
  (xin_0 => "001001100011010001", xin_1 => "001001110110111001", pass => false),
  (xin_0 => "001011010110111001", xin_1 => "000011010111111011", pass => true),
  (xin_0 => "001100100010101111", xin_1 => "001000101111100110", pass => false),
  (xin_0 => "000111001010110111", xin_1 => "000111011110111000", pass => true),
  (xin_0 => "001111010101101100", xin_1 => "001010000011000011", pass => true),
  (xin_0 => "000111110011100100", xin_1 => "001001111001110011", pass => false),
  (xin_0 => "000101001101001011", xin_1 => "001000111011111011", pass => false),
  (xin_0 => "001010101100110001", xin_1 => "000110101010101110", pass => true),
  (xin_0 => "000110010111110100", xin_1 => "000100010110100100", pass => true),
  (xin_0 => "000100101110001011", xin_1 => "001001111000001001", pass => false),
  (xin_0 => "001010101110111110", xin_1 => "000110001010001000", pass => true),
  (xin_0 => "001011100101011000", xin_1 => "000100101100001011", pass => true),
  (xin_0 => "001011100100101011", xin_1 => "000110110100011111", pass => false),
  (xin_0 => "001010010111101001", xin_1 => "001000111110011101", pass => false),
  (xin_0 => "000110010101100101", xin_1 => "000101111110100100", pass => true),
  (xin_0 => "000100111010101001", xin_1 => "001000110110010001", pass => false),
  (xin_0 => "000011111000001011", xin_1 => "000000011000111101", pass => true),
  (xin_0 => "001001100010111000", xin_1 => "000010010010111010", pass => false),
  (xin_0 => "001000001001011101", xin_1 => "000010111011011001", pass => false),
  (xin_0 => "001000101100111100", xin_1 => "000010000100011001", pass => false),
  (xin_0 => "001001101001000111", xin_1 => "000100100011011001", pass => true),
  (xin_0 => "001100010011100101", xin_1 => "001000110011010110", pass => false),
  (xin_0 => "001010010110110001", xin_1 => "000100111011011010", pass => true),
  (xin_0 => "000110000101011011", xin_1 => "000110111011100001", pass => true),
  (xin_0 => "001100101100101001", xin_1 => "000011000011100101", pass => true),
  (xin_0 => "001000000100011100", xin_1 => "000110110100010000", pass => true),
  (xin_0 => "001000101010110110", xin_1 => "000011001001010100", pass => false),
  (xin_0 => "001010100110110111", xin_1 => "000110110100111101", pass => true),
  (xin_0 => "001010100000110101", xin_1 => "001010011010111010", pass => false),
  (xin_0 => "000101110111110011", xin_1 => "001000101101100011", pass => false),
  (xin_0 => "001001100011000010", xin_1 => "000100110011000001", pass => true),
  (xin_0 => "001010001101100000", xin_1 => "000111000111111101", pass => true),
  (xin_0 => "001101010111111011", xin_1 => "000110011110110111", pass => false),
  (xin_0 => "001000000000101010", xin_1 => "000010001110001011", pass => false),
  (xin_0 => "001000101000010111", xin_1 => "000010001011101101", pass => false),
  (xin_0 => "001100111110001000", xin_1 => "000110001100000010", pass => false),
  (xin_0 => "000111100011111001", xin_1 => "000011011110100110", pass => false),
  (xin_0 => "000101011100000010", xin_1 => "001000100101110111", pass => false),
  (xin_0 => "000111001110100101", xin_1 => "001001100010110011", pass => false),
  (xin_0 => "000111010001010110", xin_1 => "000010001010101001", pass => false),
  (xin_0 => "000110100010010111", xin_1 => "000010100111100101", pass => false),
  (xin_0 => "000011100101000010", xin_1 => "000101001010100000", pass => true),
  (xin_0 => "001100010001111110", xin_1 => "000001100111000100", pass => true),
  (xin_0 => "000100111011110110", xin_1 => "000101010111100111", pass => true),
  (xin_0 => "001000110001100010", xin_1 => "000111010100001000", pass => true),
  (xin_0 => "001100010100011010", xin_1 => "000101001001001011", pass => true),
  (xin_0 => "001001000001110000", xin_1 => "000110111010111000", pass => true),
  (xin_0 => "001000110011100101", xin_1 => "000010100111110111", pass => false),
  (xin_0 => "000111100101011100", xin_1 => "000111000010100100", pass => true),
  (xin_0 => "000111101110011100", xin_1 => "001100010101111100", pass => false),
  (xin_0 => "001100100001001001", xin_1 => "000001100001011101", pass => true),
  (xin_0 => "001100001011010001", xin_1 => "001001001110111010", pass => false),
  (xin_0 => "000111111100101110", xin_1 => "000010110011001000", pass => false),
  (xin_0 => "001000000111000100", xin_1 => "000111111011101011", pass => true),
  (xin_0 => "000110001000011110", xin_1 => "000110000101011011", pass => true),
  (xin_0 => "001110011011111111", xin_1 => "001000110000110100", pass => true),
  (xin_0 => "001011011010110010", xin_1 => "001001000111011110", pass => false),
  (xin_0 => "001111110000011010", xin_1 => "001001111001000101", pass => true),
  (xin_0 => "001101000001111011", xin_1 => "001000111101101111", pass => false),
  (xin_0 => "000110000010001001", xin_1 => "000101100101100101", pass => true),
  (xin_0 => "000111001110111001", xin_1 => "000010100010010000", pass => false),
  (xin_0 => "001010100000001100", xin_1 => "001010011110110001", pass => false),
  (xin_0 => "000011111111001011", xin_1 => "000010010111100001", pass => true),
  (xin_0 => "001101011000010100", xin_1 => "000110111010111011", pass => false),
  (xin_0 => "000111000010100001", xin_1 => "001001001010010101", pass => false),
  (xin_0 => "001101010100110110", xin_1 => "000010101101111000", pass => true),
  (xin_0 => "001100011111110011", xin_1 => "000100011000011100", pass => true),
  (xin_0 => "001010101111011111", xin_1 => "000110001100101100", pass => true),
  (xin_0 => "001110100101111111", xin_1 => "001010110111101001", pass => true),
  (xin_0 => "000111100101000010", xin_1 => "000111000001110101", pass => true),
  (xin_0 => "001001000110110000", xin_1 => "001010100011000101", pass => false),
  (xin_0 => "001101110000000001", xin_1 => "000110111101000011", pass => false),
  (xin_0 => "000101100100000101", xin_1 => "000110000000010111", pass => true),
  (xin_0 => "000101010101111011", xin_1 => "000100011110011011", pass => true),
  (xin_0 => "001010011100011101", xin_1 => "001100111101001101", pass => false),
  (xin_0 => "000111101100010100", xin_1 => "000001100100011111", pass => false),
  (xin_0 => "000111111110010000", xin_1 => "000010001100000100", pass => false),
  (xin_0 => "001011000010110001", xin_1 => "001000011100101100", pass => false),
  (xin_0 => "001100011111100101", xin_1 => "000110111000110101", pass => false),
  (xin_0 => "001100100000001011", xin_1 => "000100010110111100", pass => true),
  (xin_0 => "001100110101001001", xin_1 => "000110001001010001", pass => false),
  (xin_0 => "000011010001010010", xin_1 => "000111100101001011", pass => false),
  (xin_0 => "000011011000100100", xin_1 => "000001101010001110", pass => true),
  (xin_0 => "000101000011000001", xin_1 => "000100110000010001", pass => true),
  (xin_0 => "000011110001001100", xin_1 => "000101110110011011", pass => true),
  (xin_0 => "000111000111111011", xin_1 => "000011011100110010", pass => false),
  (xin_0 => "001100111101111001", xin_1 => "001010110101100001", pass => true),
  (xin_0 => "001001111001111100", xin_1 => "000101000110100001", pass => true),
  (xin_0 => "000110110000001000", xin_1 => "000010011001111110", pass => false),
  (xin_0 => "000011001010000110", xin_1 => "000000111111000001", pass => true),
  (xin_0 => "001010001010010110", xin_1 => "000001100010011000", pass => false),
  (xin_0 => "000101011011100011", xin_1 => "000101111011110111", pass => true),
  (xin_0 => "000110011001011001", xin_1 => "001010001001001110", pass => false),
  (xin_0 => "001001000100011010", xin_1 => "000010010110001000", pass => false),
  (xin_0 => "010000000101101101", xin_1 => "001001111010100010", pass => true),
  (xin_0 => "001010000011110010", xin_1 => "000110110000100100", pass => true),
  (xin_0 => "001001010101110110", xin_1 => "000011011011001011", pass => false),
  (xin_0 => "000100100010100010", xin_1 => "000111101111010010", pass => false),
  (xin_0 => "001001101010110100", xin_1 => "000011010011101111", pass => false),
  (xin_0 => "000110111101000101", xin_1 => "000010001010111010", pass => false),
  (xin_0 => "000101010110011110", xin_1 => "000100000101001110", pass => true),
  (xin_0 => "000111011101011011", xin_1 => "001000001000000101", pass => true),
  (xin_0 => "001001001000100100", xin_1 => "000011000001101101", pass => false),
  (xin_0 => "001000000110111000", xin_1 => "001010001111111000", pass => false),
  (xin_0 => "001001011110010110", xin_1 => "000110000010010111", pass => true),
  (xin_0 => "001001101101111011", xin_1 => "000100011000111000", pass => true),
  (xin_0 => "001010111010110010", xin_1 => "000111001111110010", pass => false),
  (xin_0 => "000100110000010100", xin_1 => "000100000110001110", pass => true),
  (xin_0 => "001011110010111111", xin_1 => "000111110101111111", pass => false),
  (xin_0 => "001010101011100111", xin_1 => "000101101101000100", pass => true),
  (xin_0 => "001010001000110101", xin_1 => "000010101110111011", pass => false),
  (xin_0 => "000011011011110000", xin_1 => "000010001110100100", pass => true),
  (xin_0 => "001000011101010111", xin_1 => "000010111010101110", pass => false),
  (xin_0 => "001000111011011111", xin_1 => "000010000010101000", pass => false),
  (xin_0 => "001001100011111010", xin_1 => "000010011001101011", pass => false),
  (xin_0 => "001010110110011011", xin_1 => "001001101100100001", pass => false),
  (xin_0 => "000101010011001111", xin_1 => "000110111011010001", pass => true),
  (xin_0 => "001000111010000010", xin_1 => "000010011010000101", pass => false),
  (xin_0 => "000101010011101011", xin_1 => "000100101100101011", pass => true),
  (xin_0 => "001101010001010011", xin_1 => "001011000011010011", pass => true),
  (xin_0 => "000111011100010100", xin_1 => "001000011011110110", pass => true),
  (xin_0 => "000100011010000010", xin_1 => "000000111100100100", pass => true),
  (xin_0 => "001000100100011110", xin_1 => "001001001000001111", pass => false),
  (xin_0 => "000111001111001101", xin_1 => "000010101011000001", pass => false),
  (xin_0 => "000100010111110111", xin_1 => "000001010110010000", pass => true),
  (xin_0 => "001001111010000010", xin_1 => "001001100111000110", pass => false),
  (xin_0 => "001011110101010100", xin_1 => "000111010010010000", pass => false),
  (xin_0 => "001000011111010110", xin_1 => "000010000101100100", pass => false),
  (xin_0 => "000110111011110111", xin_1 => "000010100100010001", pass => false),
  (xin_0 => "000100100010010001", xin_1 => "000101000110111010", pass => true),
  (xin_0 => "000100101011111001", xin_1 => "001001001001010001", pass => false),
  (xin_0 => "000110010101010010", xin_1 => "001001000111111100", pass => false),
  (xin_0 => "001100001001101111", xin_1 => "000101000111110101", pass => true),
  (xin_0 => "000110111011010101", xin_1 => "000101001000101100", pass => true),
  (xin_0 => "001000101110010111", xin_1 => "000010001000000011", pass => false),
  (xin_0 => "001011111000110011", xin_1 => "000111011011101110", pass => false),
  (xin_0 => "001101010010111001", xin_1 => "001000001010011011", pass => false),
  (xin_0 => "001000110010011011", xin_1 => "000001101010100011", pass => false),
  (xin_0 => "001001001011001001", xin_1 => "000010010110111101", pass => false),
  (xin_0 => "001000110010011111", xin_1 => "000001111100110101", pass => false),
  (xin_0 => "001001100101001010", xin_1 => "000011010011100010", pass => false),
  (xin_0 => "000100110010011000", xin_1 => "000101100010110000", pass => true),
  (xin_0 => "000111110010101110", xin_1 => "000010101011100010", pass => false),
  (xin_0 => "000111010011110111", xin_1 => "000010101111111010", pass => false),
  (xin_0 => "001000011001011110", xin_1 => "001000101000011010", pass => true),
  (xin_0 => "001010001001100111", xin_1 => "000111101010101000", pass => true),
  (xin_0 => "001011000101100010", xin_1 => "001011001101100110", pass => false),
  (xin_0 => "001001011100001111", xin_1 => "000010111111110100", pass => false),
  (xin_0 => "001010000111101000", xin_1 => "000101000010101001", pass => true),
  (xin_0 => "001100001100100100", xin_1 => "001001101100010110", pass => false),
  (xin_0 => "000011111010000110", xin_1 => "000100101001010011", pass => true),
  (xin_0 => "001000110100111101", xin_1 => "000100111000100111", pass => true),
  (xin_0 => "000100110100011110", xin_1 => "001010000000110011", pass => false),
  (xin_0 => "001011000111100011", xin_1 => "000011000010111000", pass => true),
  (xin_0 => "001011110001011010", xin_1 => "001000001101101010", pass => false),
  (xin_0 => "000100110111100111", xin_1 => "001000111100100011", pass => false),
  (xin_0 => "000111011001111111", xin_1 => "001001101111000001", pass => false),
  (xin_0 => "001100001101011100", xin_1 => "000111000111101000", pass => false),
  (xin_0 => "001101010110110110", xin_1 => "000111001011111011", pass => false),
  (xin_0 => "000110010101011111", xin_1 => "000110100010001101", pass => true),
  (xin_0 => "001010110011000100", xin_1 => "001010000001100111", pass => false),
  (xin_0 => "001011011000011011", xin_1 => "001000000011111010", pass => false),
  (xin_0 => "001010110000011001", xin_1 => "000100100100010000", pass => true),
  (xin_0 => "001010001011011000", xin_1 => "001011100000100000", pass => false),
  (xin_0 => "001100100000011110", xin_1 => "000010100101100010", pass => true),
  (xin_0 => "001010001010010010", xin_1 => "000010010100101100", pass => false),
  (xin_0 => "000110111110000010", xin_1 => "001001001111000010", pass => false),
  (xin_0 => "001010001110011101", xin_1 => "000010111010011000", pass => false),
  (xin_0 => "001011011011011011", xin_1 => "001001101110000111", pass => false),
  (xin_0 => "001001001010101000", xin_1 => "000101101111000010", pass => true),
  (xin_0 => "000110111001111110", xin_1 => "000101000100111110", pass => true),
  (xin_0 => "000111011001011100", xin_1 => "000101100011001000", pass => true),
  (xin_0 => "001001100001110101", xin_1 => "000011100111001010", pass => false),
  (xin_0 => "000110110011111001", xin_1 => "000110000001101110", pass => true),
  (xin_0 => "000110110011000001", xin_1 => "000110110100110010", pass => true),
  (xin_0 => "000100001111011100", xin_1 => "000111000111100100", pass => false),
  (xin_0 => "001000101000110111", xin_1 => "000011100010100001", pass => false),
  (xin_0 => "001011111001001011", xin_1 => "000011000001100110", pass => true),
  (xin_0 => "001011101000011010", xin_1 => "001000110110000000", pass => false),
  (xin_0 => "001100011001111101", xin_1 => "000010011011111001", pass => true),
  (xin_0 => "001001111011001101", xin_1 => "001001101110100101", pass => false),
  (xin_0 => "000111110101010110", xin_1 => "001010110010111000", pass => false),
  (xin_0 => "000101110100000111", xin_1 => "000010010001111001", pass => false),
  (xin_0 => "001000001010000001", xin_1 => "000001010110100110", pass => false),
  (xin_0 => "000100100101011001", xin_1 => "000101010111000111", pass => true),
  (xin_0 => "001011001011010110", xin_1 => "000011011100000100", pass => true),
  (xin_0 => "010000011101100010", xin_1 => "001001110000001110", pass => true),
  (xin_0 => "000011111011101110", xin_1 => "000010001101010110", pass => true),
  (xin_0 => "001101101101110110", xin_1 => "000101110001000010", pass => false),
  (xin_0 => "001100001011101010", xin_1 => "000111010111011111", pass => false),
  (xin_0 => "001011111010000111", xin_1 => "000100010101000011", pass => true),
  (xin_0 => "001111101111100100", xin_1 => "001011001101010110", pass => true),
  (xin_0 => "000101011100111101", xin_1 => "000100111110111111", pass => true),
  (xin_0 => "001110001011000000", xin_1 => "000011110000110001", pass => false),
  (xin_0 => "000110111010010001", xin_1 => "000110100111101101", pass => true),
  (xin_0 => "001000111001100011", xin_1 => "000001100001110111", pass => false),
  (xin_0 => "001100011001000010", xin_1 => "001001010000100101", pass => false),
  (xin_0 => "000100011001000011", xin_1 => "001001000101110111", pass => false),
  (xin_0 => "001000000011100001", xin_1 => "001010100111110110", pass => false),
  (xin_0 => "000111000110100111", xin_1 => "000011001001100110", pass => false),
  (xin_0 => "001000011101100000", xin_1 => "000101001011010001", pass => true),
  (xin_0 => "001100110010110101", xin_1 => "000100110000000000", pass => true),
  (xin_0 => "000101111001100011", xin_1 => "000101000000101111", pass => true),
  (xin_0 => "000110000011110010", xin_1 => "001000111110110010", pass => false),
  (xin_0 => "001110000100010011", xin_1 => "001010010001010110", pass => true),
  (xin_0 => "001011011011111011", xin_1 => "001000111000110101", pass => false),
  (xin_0 => "000011100111111100", xin_1 => "000101010111010110", pass => true),
  (xin_0 => "000100101001010111", xin_1 => "001000011111010001", pass => false),
  (xin_0 => "001000010000101011", xin_1 => "000011101001101000", pass => false),
  (xin_0 => "000100100100000100", xin_1 => "000011111000111101", pass => true),
  (xin_0 => "001000001101011111", xin_1 => "000101111000001011", pass => true),
  (xin_0 => "000011101111101111", xin_1 => "000010011001111101", pass => true),
  (xin_0 => "001000010101000110", xin_1 => "000101100100011100", pass => true),
  (xin_0 => "001101111010111110", xin_1 => "000101010110011000", pass => false),
  (xin_0 => "000100110100010010", xin_1 => "000110100000010010", pass => true),
  (xin_0 => "001000101001100010", xin_1 => "000100111000011111", pass => true),
  (xin_0 => "000111111100111011", xin_1 => "000001101011000010", pass => false),
  (xin_0 => "000110010000111110", xin_1 => "001010111011111100", pass => false),
  (xin_0 => "000011010001100010", xin_1 => "000010111011010000", pass => true),
  (xin_0 => "001100101111001111", xin_1 => "001001000100100100", pass => false),
  (xin_0 => "000101111100011000", xin_1 => "000110000111100100", pass => true),
  (xin_0 => "001001010000100010", xin_1 => "000101100110001001", pass => true),
  (xin_0 => "001010101101101011", xin_1 => "000010101000101001", pass => true),
  (xin_0 => "001000000010100100", xin_1 => "000010010001100101", pass => false),
  (xin_0 => "010000100111000111", xin_1 => "001001101101010001", pass => true),
  (xin_0 => "000110000100101000", xin_1 => "000110110011110100", pass => true),
  (xin_0 => "001100010101000011", xin_1 => "000010110111100111", pass => true),
  (xin_0 => "001000110011000100", xin_1 => "001011000101011101", pass => false),
  (xin_0 => "001010111100000100", xin_1 => "001011010111100001", pass => false),
  (xin_0 => "000100011000101001", xin_1 => "000101001010001000", pass => true),
  (xin_0 => "000111010000110110", xin_1 => "000010001000011100", pass => false),
  (xin_0 => "001000111001111111", xin_1 => "000010111101100011", pass => false),
  (xin_0 => "001100110101110101", xin_1 => "000100010011101010", pass => true),
  (xin_0 => "001011100001101101", xin_1 => "001000101101011101", pass => false),
  (xin_0 => "001010000010010001", xin_1 => "000010101011010001", pass => false),
  (xin_0 => "001010000101010110", xin_1 => "000010100100100010", pass => false),
  (xin_0 => "001011001010100001", xin_1 => "001001101110100001", pass => false),
  (xin_0 => "000101001100110111", xin_1 => "000101100001110010", pass => true),
  (xin_0 => "001011110110001111", xin_1 => "000010110100010011", pass => true),
  (xin_0 => "001011110100110001", xin_1 => "001000000010001000", pass => false),
  (xin_0 => "001001010111110101", xin_1 => "000100111101111001", pass => true),
  (xin_0 => "000010110010110111", xin_1 => "001000010010011110", pass => false),
  (xin_0 => "000110101111001011", xin_1 => "000010110001110111", pass => false),
  (xin_0 => "001001111111111000", xin_1 => "001001000011101110", pass => false),
  (xin_0 => "001101110011110011", xin_1 => "000101010101100000", pass => false),
  (xin_0 => "001000100011011001", xin_1 => "000011000110011001", pass => false),
  (xin_0 => "001010000100000111", xin_1 => "000011101110010110", pass => true),
  (xin_0 => "000110111010011000", xin_1 => "000011110010100110", pass => false),
  (xin_0 => "001110001001011010", xin_1 => "001010110010100001", pass => true),
  (xin_0 => "001011011111100100", xin_1 => "000110101101110100", pass => false),
  (xin_0 => "001100011111001101", xin_1 => "001010010100011000", pass => false),
  (xin_0 => "001011010010110011", xin_1 => "000011101100110100", pass => true),
  (xin_0 => "001100100000100110", xin_1 => "000110001100111010", pass => false),
  (xin_0 => "001000100101000000", xin_1 => "000001000101011001", pass => false),
  (xin_0 => "000110010110101000", xin_1 => "000011000011101101", pass => false),
  (xin_0 => "001001101011010011", xin_1 => "000010111000110011", pass => false),
  (xin_0 => "001000111001010000", xin_1 => "000010011000101001", pass => false),
  (xin_0 => "001110010100000111", xin_1 => "000100100001111111", pass => false),
  (xin_0 => "000111000100010010", xin_1 => "000101111010011101", pass => true),
  (xin_0 => "001100011111110110", xin_1 => "000101101111101110", pass => false),
  (xin_0 => "000110101100011100", xin_1 => "000100111010111100", pass => true),
  (xin_0 => "001001001110111111", xin_1 => "000100011011001110", pass => true),
  (xin_0 => "000101001101110100", xin_1 => "000111110010000001", pass => false),
  (xin_0 => "001000000011011011", xin_1 => "000010111111010101", pass => false),
  (xin_0 => "000101000101110001", xin_1 => "000110000101101011", pass => true),
  (xin_0 => "000111001100100111", xin_1 => "000100100100010101", pass => true),
  (xin_0 => "000101101010101110", xin_1 => "001001010011110110", pass => false),
  (xin_0 => "000110010011011111", xin_1 => "000100101000111011", pass => true),
  (xin_0 => "001100101001001000", xin_1 => "000110011110111100", pass => false),
  (xin_0 => "000111011101011000", xin_1 => "000011011100100000", pass => false),
  (xin_0 => "000111110011011000", xin_1 => "001010001110011010", pass => false),
  (xin_0 => "000100011101001101", xin_1 => "000001110000110110", pass => true),
  (xin_0 => "001000100110001101", xin_1 => "000010111110110011", pass => false),
  (xin_0 => "001000001100110111", xin_1 => "001010010111110101", pass => false),
  (xin_0 => "001110100110010111", xin_1 => "001001100010000001", pass => true),
  (xin_0 => "001010111011000011", xin_1 => "001000010111001110", pass => false),
  (xin_0 => "000101001001001000", xin_1 => "001001101000010000", pass => false),
  (xin_0 => "001010100010001010", xin_1 => "001010000111001101", pass => false),
  (xin_0 => "001001000010011010", xin_1 => "000010110101001110", pass => false),
  (xin_0 => "001010010100010011", xin_1 => "001010011101101110", pass => false),
  (xin_0 => "001001101011100000", xin_1 => "000110101111110111", pass => true),
  (xin_0 => "000101110010010000", xin_1 => "000100110100100011", pass => true),
  (xin_0 => "000111101010000010", xin_1 => "000011001011001001", pass => false),
  (xin_0 => "001001000110000001", xin_1 => "000101000010110100", pass => true),
  (xin_0 => "001000110101101001", xin_1 => "000010111010111111", pass => false),
  (xin_0 => "000111110101111110", xin_1 => "001000010001000111", pass => true),
  (xin_0 => "001100100100100001", xin_1 => "000110001110000011", pass => false),
  (xin_0 => "000111010001001101", xin_1 => "001010010110110101", pass => false),
  (xin_0 => "000100000011100110", xin_1 => "000110000101100101", pass => true),
  (xin_0 => "001110001111110010", xin_1 => "000111100110100000", pass => false),
  (xin_0 => "000111001000011100", xin_1 => "000101110111101011", pass => true),
  (xin_0 => "000011101010110001", xin_1 => "001000111010101111", pass => false),
  (xin_0 => "001001010001001111", xin_1 => "000100101000111100", pass => true),
  (xin_0 => "000101101101111000", xin_1 => "000110101100100000", pass => true),
  (xin_0 => "001100100001110101", xin_1 => "000111100111101100", pass => false),
  (xin_0 => "001001011011000001", xin_1 => "000011110100100110", pass => false),
  (xin_0 => "001000100010000001", xin_1 => "000011100101100001", pass => false),
  (xin_0 => "001000111111011100", xin_1 => "000011010010001001", pass => false),
  (xin_0 => "001110001000001111", xin_1 => "000101111010110011", pass => false),
  (xin_0 => "001010001001000111", xin_1 => "001001010011100001", pass => false),
  (xin_0 => "001011000111110010", xin_1 => "000100100001111011", pass => true),
  (xin_0 => "000110101001101000", xin_1 => "000111000100010100", pass => true),
  (xin_0 => "000100111100011111", xin_1 => "000011101101111000", pass => true),
  (xin_0 => "000101000011111011", xin_1 => "000101010010010011", pass => true),
  (xin_0 => "000100110000011010", xin_1 => "000010110000001011", pass => true),
  (xin_0 => "001011111011101010", xin_1 => "000111111001000110", pass => false),
  (xin_0 => "001100011010110011", xin_1 => "000111010100110000", pass => false),
  (xin_0 => "001010101010111000", xin_1 => "001001001011111000", pass => false),
  (xin_0 => "001001011011010011", xin_1 => "000010110010110110", pass => false),
  (xin_0 => "000100011001110100", xin_1 => "000011111000010010", pass => true),
  (xin_0 => "000111101101001000", xin_1 => "000101001011001111", pass => true),
  (xin_0 => "001010101110101111", xin_1 => "000101100101100011", pass => true),
  (xin_0 => "000110011110010010", xin_1 => "000100001101010011", pass => true),
  (xin_0 => "001000010001001101", xin_1 => "000001100010000000", pass => false),
  (xin_0 => "000100100100010111", xin_1 => "000100010100101101", pass => true),
  (xin_0 => "000011110110100010", xin_1 => "000100010011101001", pass => true),
  (xin_0 => "000100001010000100", xin_1 => "000001100110000010", pass => true),
  (xin_0 => "000110110001101000", xin_1 => "000101010000100101", pass => true),
  (xin_0 => "000110001111101110", xin_1 => "000001011011000100", pass => false),
  (xin_0 => "001000111000011100", xin_1 => "000101110011001001", pass => true),
  (xin_0 => "000111011100001001", xin_1 => "000010001010001000", pass => false),
  (xin_0 => "001011000001011010", xin_1 => "000010100110011010", pass => true),
  (xin_0 => "001011010110010001", xin_1 => "001000011111010110", pass => false),
  (xin_0 => "001001110110000010", xin_1 => "001001000100001001", pass => false),
  (xin_0 => "001011001110101010", xin_1 => "000100011001101110", pass => true),
  (xin_0 => "001101111010110011", xin_1 => "000101100010110111", pass => false),
  (xin_0 => "001110011100010010", xin_1 => "000101011111010111", pass => false),
  (xin_0 => "000111010101000010", xin_1 => "000111101010101010", pass => true),
  (xin_0 => "000101000001001101", xin_1 => "000011101001100001", pass => true),
  (xin_0 => "001000010011000011", xin_1 => "000011000000101001", pass => false),
  (xin_0 => "000110001100101001", xin_1 => "000010010001011100", pass => false),
  (xin_0 => "000111000100001100", xin_1 => "000100100111110001", pass => true),
  (xin_0 => "001001100110010000", xin_1 => "000110111000001100", pass => true),
  (xin_0 => "000110000011101101", xin_1 => "001001110111110001", pass => false),
  (xin_0 => "000100100000001010", xin_1 => "000100011010001111", pass => true),
  (xin_0 => "001000010000010011", xin_1 => "000101000101110010", pass => true),
  (xin_0 => "001000010101111111", xin_1 => "000110100100000000", pass => true),
  (xin_0 => "001000010000111000", xin_1 => "000001101100010100", pass => false),
  (xin_0 => "001100000000001010", xin_1 => "001000010110110110", pass => false),
  (xin_0 => "000110111101111011", xin_1 => "001000011100000101", pass => true),
  (xin_0 => "001000110101111100", xin_1 => "000011110100110000", pass => false),
  (xin_0 => "001000001101000000", xin_1 => "000111101110111110", pass => true),
  (xin_0 => "001100011101110000", xin_1 => "001000100000111100", pass => false),
  (xin_0 => "000100011100110110", xin_1 => "000110100110000001", pass => true),
  (xin_0 => "000111010110001010", xin_1 => "000011001000101110", pass => false),
  (xin_0 => "001000110110101100", xin_1 => "000010111111000001", pass => false),
  (xin_0 => "000111101011010101", xin_1 => "000010010001110110", pass => false),
  (xin_0 => "001011010001101110", xin_1 => "001001111010001000", pass => false),
  (xin_0 => "000101100011000011", xin_1 => "001000010101010001", pass => false),
  (xin_0 => "000111011000111110", xin_1 => "001010011111111111", pass => false),
  (xin_0 => "001100001100000001", xin_1 => "000111010111100110", pass => false),
  (xin_0 => "000101110110010011", xin_1 => "000110000110111110", pass => true),
  (xin_0 => "001001001011111001", xin_1 => "000010101111001111", pass => false),
  (xin_0 => "000011011000000101", xin_1 => "000010101010000111", pass => true),
  (xin_0 => "001010100100111100", xin_1 => "001001110011110111", pass => false),
  (xin_0 => "001000011110111011", xin_1 => "000010011101011011", pass => false),
  (xin_0 => "001001101011000110", xin_1 => "000100110110111011", pass => true),
  (xin_0 => "000110111011011101", xin_1 => "000110001110011101", pass => true),
  (xin_0 => "001101010011110001", xin_1 => "001010110010010101", pass => true),
  (xin_0 => "001000011100010000", xin_1 => "000010110101011001", pass => false),
  (xin_0 => "000101101001000110", xin_1 => "000101011110111111", pass => true),
  (xin_0 => "001100000000101000", xin_1 => "001000111101011011", pass => false),
  (xin_0 => "001011100000000011", xin_1 => "001001010111000111", pass => false),
  (xin_0 => "001010110101100100", xin_1 => "001011111001010110", pass => false),
  (xin_0 => "000111111011111110", xin_1 => "000011001011011011", pass => false),
  (xin_0 => "001110110001010010", xin_1 => "000100000111010010", pass => false),
  (xin_0 => "001100010000111001", xin_1 => "000101111110011100", pass => false),
  (xin_0 => "000011110011011010", xin_1 => "000011101010100011", pass => true),
  (xin_0 => "001010111111100011", xin_1 => "000011011110010110", pass => true),
  (xin_0 => "000101100101100110", xin_1 => "000111101001111000", pass => true),
  (xin_0 => "000100011011011110", xin_1 => "000011000010010100", pass => true),
  (xin_0 => "001111010000110011", xin_1 => "001001101001111010", pass => true),
  (xin_0 => "000111111000000001", xin_1 => "000010000001001111", pass => false),
  (xin_0 => "000110101110011000", xin_1 => "001010010101111001", pass => false),
  (xin_0 => "001000001110010101", xin_1 => "001000000111110001", pass => true),
  (xin_0 => "001100000101010101", xin_1 => "000000111001000100", pass => true),
  (xin_0 => "001000111001000001", xin_1 => "001000010111011100", pass => true),
  (xin_0 => "000100111100111001", xin_1 => "000010111011101111", pass => true),
  (xin_0 => "001000011011100111", xin_1 => "000100010010001001", pass => false),
  (xin_0 => "001100110110001111", xin_1 => "001000111001011001", pass => false),
  (xin_0 => "001000100000100110", xin_1 => "000010100000100100", pass => false),
  (xin_0 => "001001100101010001", xin_1 => "000010100011010101", pass => false),
  (xin_0 => "000111000100010111", xin_1 => "000111010110010110", pass => true),
  (xin_0 => "001011111000110010", xin_1 => "000011011000101111", pass => true),
  (xin_0 => "001001001000000110", xin_1 => "000010011000111110", pass => false),
  (xin_0 => "001011100110010000", xin_1 => "000101000101110000", pass => true),
  (xin_0 => "000110101000011110", xin_1 => "000101011111111000", pass => true),
  (xin_0 => "000111111110100010", xin_1 => "001011010001100000", pass => false),
  (xin_0 => "000110110100111011", xin_1 => "001010000001111100", pass => false),
  (xin_0 => "001000111000100001", xin_1 => "000010010101101000", pass => false),
  (xin_0 => "001011001110011010", xin_1 => "001001001011101110", pass => false),
  (xin_0 => "001000101101110100", xin_1 => "001011001100110111", pass => false),
  (xin_0 => "001000011000110110", xin_1 => "001010001101010010", pass => false),
  (xin_0 => "001000010101001111", xin_1 => "000101100000111001", pass => true),
  (xin_0 => "001000010111111111", xin_1 => "000011000111001101", pass => false),
  (xin_0 => "000111110101111111", xin_1 => "000011000011101000", pass => false),
  (xin_0 => "001010001100110001", xin_1 => "000100001111010001", pass => true),
  (xin_0 => "001010100111101111", xin_1 => "000011000010101111", pass => true),
  (xin_0 => "000111011110110001", xin_1 => "001010101110000101", pass => false),
  (xin_0 => "001100001010100011", xin_1 => "000110010111111100", pass => false),
  (xin_0 => "000011110110010111", xin_1 => "000001011010100000", pass => true),
  (xin_0 => "000110001000101001", xin_1 => "000110100011011110", pass => true),
  (xin_0 => "001100100111001001", xin_1 => "000100100010111101", pass => true),
  (xin_0 => "001000111101100011", xin_1 => "000101110110001011", pass => true),
  (xin_0 => "000111110011111110", xin_1 => "001010011100110010", pass => false),
  (xin_0 => "000111110000011111", xin_1 => "001001110011001001", pass => false),
  (xin_0 => "000110010000000111", xin_1 => "000010101111001100", pass => false),
  (xin_0 => "000111000110011001", xin_1 => "000011010111110111", pass => false),
  (xin_0 => "001000110000110110", xin_1 => "000001011100011100", pass => false),
  (xin_0 => "001010101111010100", xin_1 => "000010111110001111", pass => true),
  (xin_0 => "000010001110100010", xin_1 => "000110011111010100", pass => false),
  (xin_0 => "001010001100111011", xin_1 => "000001110010100110", pass => false),
  (xin_0 => "001010100010011011", xin_1 => "001001101110001100", pass => false),
  (xin_0 => "001001011001101000", xin_1 => "000100001111100100", pass => true),
  (xin_0 => "001100100011011111", xin_1 => "000111111010011011", pass => false),
  (xin_0 => "001001110010001110", xin_1 => "000001110100111011", pass => false),
  (xin_0 => "000111000110001001", xin_1 => "000111110010111010", pass => true),
  (xin_0 => "001000110010111110", xin_1 => "000010010000000001", pass => false),
  (xin_0 => "001010010101011001", xin_1 => "001000101000011111", pass => false),
  (xin_0 => "000110100010001001", xin_1 => "000011000000010011", pass => false),
  (xin_0 => "000110011110100010", xin_1 => "000011000010000010", pass => false),
  (xin_0 => "001000110111110010", xin_1 => "000101001111101010", pass => true),
  (xin_0 => "000011100000001100", xin_1 => "000010011001010100", pass => true),
  (xin_0 => "001111000110010010", xin_1 => "001001100100100110", pass => true),
  (xin_0 => "000101000110000111", xin_1 => "000101011000110110", pass => true),
  (xin_0 => "001001000100111100", xin_1 => "000011000011101010", pass => false),
  (xin_0 => "001100101111001010", xin_1 => "001011001010001010", pass => true),
  (xin_0 => "000110111111010001", xin_1 => "000010001100110100", pass => false),
  (xin_0 => "001101000010100110", xin_1 => "000110100000001101", pass => false),
  (xin_0 => "000100111001101101", xin_1 => "001001110110111001", pass => false),
  (xin_0 => "000111100010101111", xin_1 => "000011110011011011", pass => false),
  (xin_0 => "001100001111000011", xin_1 => "001001011101110010", pass => false),
  (xin_0 => "000111000001000010", xin_1 => "000010110010001010", pass => false),
  (xin_0 => "000111011011000101", xin_1 => "000111001000001110", pass => true),
  (xin_0 => "001010001011100001", xin_1 => "000101001101100010", pass => true),
  (xin_0 => "000101100011001011", xin_1 => "000110100110111111", pass => true),
  (xin_0 => "000100110001010100", xin_1 => "000100111010111000", pass => true),
  (xin_0 => "000110011111111111", xin_1 => "000011100101001001", pass => false),
  (xin_0 => "001101111001010110", xin_1 => "000111111101001110", pass => false),
  (xin_0 => "001001101111011000", xin_1 => "000001010111010010", pass => false),
  (xin_0 => "001010000100010011", xin_1 => "000101010001011011", pass => true),
  (xin_0 => "000111111111111011", xin_1 => "000011010100110011", pass => false),
  (xin_0 => "000111011110100111", xin_1 => "000011101110001011", pass => false),
  (xin_0 => "000111001110100101", xin_1 => "001000001000001000", pass => true),
  (xin_0 => "001010011011100101", xin_1 => "000010101111100011", pass => false),
  (xin_0 => "001000011100000011", xin_1 => "000100100011011101", pass => true),
  (xin_0 => "001011111101101100", xin_1 => "000010110010100001", pass => true),
  (xin_0 => "001000011011011011", xin_1 => "000010111000100010", pass => false),
  (xin_0 => "000111100010011011", xin_1 => "000100100000011111", pass => true),
  (xin_0 => "001011111100111000", xin_1 => "000011110001111001", pass => true),
  (xin_0 => "001001011111101100", xin_1 => "000011000111100100", pass => false),
  (xin_0 => "000010111110111011", xin_1 => "000111011010110001", pass => false),
  (xin_0 => "001010111100110001", xin_1 => "000101101010001011", pass => true),
  (xin_0 => "001010000110010001", xin_1 => "000011000100111000", pass => false),
  (xin_0 => "001100011101011100", xin_1 => "000111001010001011", pass => false),
  (xin_0 => "000111000100110001", xin_1 => "000100010011110001", pass => false),
  (xin_0 => "000101111000011000", xin_1 => "000011011000010101", pass => false),
  (xin_0 => "000111100011011001", xin_1 => "001001101111011101", pass => false),
  (xin_0 => "000111111110100101", xin_1 => "000111111011011001", pass => true),
  (xin_0 => "001001000111111000", xin_1 => "000101110100101000", pass => true),
  (xin_0 => "001111110001110010", xin_1 => "001010110010100011", pass => true),
  (xin_0 => "001100010011101001", xin_1 => "000100110101011100", pass => true),
  (xin_0 => "001000011001111010", xin_1 => "000010011101111110", pass => false),
  (xin_0 => "001011011011011100", xin_1 => "000100100110000000", pass => true),
  (xin_0 => "001100010001111001", xin_1 => "000010110001010111", pass => true),
  (xin_0 => "001001001110111011", xin_1 => "000010111111100010", pass => false),
  (xin_0 => "001011001100011101", xin_1 => "001000000110100011", pass => false),
  (xin_0 => "001011010110101100", xin_1 => "001010111101110010", pass => false),
  (xin_0 => "001100010111001010", xin_1 => "000111110001000111", pass => false),
  (xin_0 => "001010100101011000", xin_1 => "001000001111000100", pass => false),
  (xin_0 => "001001100011011011", xin_1 => "000110010100011110", pass => true),
  (xin_0 => "001100010001101111", xin_1 => "000011001010011100", pass => true),
  (xin_0 => "001011001010010111", xin_1 => "000111010001011010", pass => false),
  (xin_0 => "001000101111110110", xin_1 => "001011001011100010", pass => false),
  (xin_0 => "000101011110111011", xin_1 => "001010100101101001", pass => false),
  (xin_0 => "001101101011100010", xin_1 => "000100100001101011", pass => false),
  (xin_0 => "000110001011000001", xin_1 => "001010010011110000", pass => false),
  (xin_0 => "000110100000011001", xin_1 => "000110001110000100", pass => true),
  (xin_0 => "000101010101010110", xin_1 => "000011011111111110", pass => true),
  (xin_0 => "000110011111100100", xin_1 => "000101101010001001", pass => true),
  (xin_0 => "000011010011110010", xin_1 => "001000000110000011", pass => false),
  (xin_0 => "001011110101010111", xin_1 => "000110011100110110", pass => false),
  (xin_0 => "001001001101011100", xin_1 => "000011101010010011", pass => false),
  (xin_0 => "000111011101010001", xin_1 => "001010101001101100", pass => false),
  (xin_0 => "001110001110110100", xin_1 => "000100010001011101", pass => false),
  (xin_0 => "001001101000010001", xin_1 => "000101011001000111", pass => true),
  (xin_0 => "001001000101001000", xin_1 => "000111110110111001", pass => true),
  (xin_0 => "001001110111001110", xin_1 => "001011110100100111", pass => false),
  (xin_0 => "000100001011110010", xin_1 => "000110000001000110", pass => true),
  (xin_0 => "001100000000010010", xin_1 => "111111111010010001", pass => true),
  (xin_0 => "000111011110010001", xin_1 => "001010111000010101", pass => false),
  (xin_0 => "000110011110111011", xin_1 => "000101010100100000", pass => true),
  (xin_0 => "000111000010100010", xin_1 => "001010100000101001", pass => false),
  (xin_0 => "000100100110110001", xin_1 => "000101000010101111", pass => true),
  (xin_0 => "000110010110110110", xin_1 => "000110110110111000", pass => true),
  (xin_0 => "001001111111100100", xin_1 => "001010110101011001", pass => false),
  (xin_0 => "001011001001110001", xin_1 => "000110010100111100", pass => true),
  (xin_0 => "001001101111011101", xin_1 => "001000101100110100", pass => false),
  (xin_0 => "001001011110000000", xin_1 => "000010011110000111", pass => false),
  (xin_0 => "001000000101001000", xin_1 => "001011011000001110", pass => false),
  (xin_0 => "001111001010000110", xin_1 => "000100110110010111", pass => false),
  (xin_0 => "001010010000000001", xin_1 => "001000011000101011", pass => false),
  (xin_0 => "000111110000000100", xin_1 => "001010101111010001", pass => false),
  (xin_0 => "000110010011011110", xin_1 => "000111001100001011", pass => true),
  (xin_0 => "001101000001111110", xin_1 => "001000101111111111", pass => false),
  (xin_0 => "001001011000001011", xin_1 => "000101110001000111", pass => true),
  (xin_0 => "001100001011101011", xin_1 => "000010111000000001", pass => true),
  (xin_0 => "001001110101001101", xin_1 => "000011010111101001", pass => false),
  (xin_0 => "001001101101011100", xin_1 => "000110111000001110", pass => true),
  (xin_0 => "000111010001001101", xin_1 => "000111111111110001", pass => true),
  (xin_0 => "000110100101001010", xin_1 => "001010000010110111", pass => false),
  (xin_0 => "000110111000000101", xin_1 => "000011000110110111", pass => false),
  (xin_0 => "001000100000111010", xin_1 => "000010110110000000", pass => false),
  (xin_0 => "000101010000000111", xin_1 => "000010110100000011", pass => true),
  (xin_0 => "000110110010010111", xin_1 => "000100011111101001", pass => true),
  (xin_0 => "000110101000000001", xin_1 => "000100000101011000", pass => false)
);
  signal clk : std_logic := '0';
  signal rst : std_logic := '1';
  signal rst1 : std_logic := '1';
  signal rst2 : std_logic := '0';
  signal ready : std_logic;
  signal done : std_logic;

  signal result_sign : std_logic ;
  signal xin_input : signed(XIN_DATA_BITS -1 downto 0):= (others=>'0');
  signal xin_addr  :  unsigned(XIN_ADDR_BITS-1 downto 0);

  signal xin_0 : signed(XIN_DATA_BITS -1 downto 0):= (others=>'0');
  signal xin_1 : signed(XIN_DATA_BITS -1 downto 0):= (others=>'0');
  signal errors: integer := 0;
  signal pass : boolean;
  signal do_rst: boolean := true;

  component csvm is
    port(
        clk         : in std_logic;
        rst         : in std_logic;
	xin  : in signed(XIN_DATA_BITS -1 downto 0);
	xin_addr    : out unsigned(XIN_ADDR_BITS-1 downto 0);
        ready       : out std_logic;
	valid_answer: out std_logic;

        result_sign : out std_logic
  );

  end component csvm;
  
begin  

  CSVM_COMP: csvm
    port map (
        clk    => clk,
        rst    => rst,
        xin   =>xin_input,
	xin_addr    => xin_addr,--: out unsigned(XIN_ADDR_BITS-1 downto 0);
        ready  => ready,
        valid_answer => done,
        result_sign => result_sign
    );
  clk  <= not clk after 5 ns;
  rst  <= rst1 or rst2;
  rst1 <= '0' after 20 ns;
  rst2 <= done;

  --process(do_reset)
  --begin
    
  --end process;

  verify: process
    variable vector: test_vector;
    variable errors: integer := 0;
  begin
    for i in test_vectors'range loop
      vector := test_vectors(i);
      xin_0 <= vector.xin_0;
      xin_1 <= vector.xin_1;
      pass <= vector.pass;
      wait until (done'event and done = '1');
    end loop;
  end process verify;

  process(xin_addr,xin_0,xin_1)
  begin
    if( xin_addr = "0") then
      --xin_input <= "001011011100110110";  --0
      --xin_input <=  "001011110001011010" ; --3
      xin_input <= xin_0;
      --                  1011011100110110
    else
      --xin_input <= "000010011110001111";  --0
      --xin_input <=  "000111100111011000"; --3
      xin_input <= xin_1;
    end if;
  end process;

  process(done)
    variable OLine : Line;
  begin
    if(done = '1') then
      if(result_sign = '1') then
        write(OLine, string'("minus"));
        writeline(output, OLine);
      else
        write(OLine, string'("plus"));
        writeline(output, OLine);

      end if;
      --assert FALSE --stop simulation
      --  report "FInished!" severity NOTE;
      assert(result_sign = '1' and pass = false)
        report "Sign mismatch: result_sign is positive, should be negative";
      assert(result_sign = '0' and pass = true)
        report "Sign mismatch: result_sign is negative, should be positive";

    end if;
    
  end process;
 

end testbench;








